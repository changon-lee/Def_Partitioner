module aes_aes_die_15 ( n1, n11, n1109, n1114, n1212, n1213, n1215, n1216, n1219, 
       n1220, n1221, n129, n13, n131, n133, n135, n137, n139, 
       n141, n143, n145, n147, n149, n15, n151, n153, n155, 
       n157, n159, n161, n163, n165, n167, n169, n17, n171, 
       n173, n175, n177, n179, n181, n183, n185, n187, n189, 
       n19, n191, n21, n23, n25, n27, n29, n3, n31, 
       n33, n35, n37, n39, n41, n43, n45, n47, n49, 
       n5, n51, n53, n55, n57, n59, n61, n63, n7, 
       n9, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, 
       sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa11_sr_0, 
       sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa13_sr_0, sa13_sr_1, 
       sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, 
       sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, 
       sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, 
       sa31_sr_5, sa31_sr_6, sa31_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, 
       sa33_sr_6, sa33_sr_7, u0_n13, u0_n250, u0_n254, u0_n258, u0_n264, u0_n33, u0_n35, 
       u0_n37, u0_n39, u0_n43, u0_n7, w1_0, w1_1, w1_10, w1_11, w1_12, 
       w1_13, w1_14, w1_15, w1_16, w1_17, w1_18, w1_19, w1_2, w1_20, 
       w1_21, w1_22, w1_23, w1_24, w1_25, w1_26, w1_27, w1_28, w1_29, 
       w1_3, w1_30, w1_31, w1_4, w1_5, w1_6, w1_7, w1_8, w1_9, 
       w2_10, w2_12, w2_13, w2_14, w2_15, w2_25, w2_28, w3_0, w3_1, 
       w3_10, w3_11, w3_16, w3_17, w3_18, w3_19, w3_2, w3_20, w3_21, 
       w3_22, w3_23, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, w3_3, 
       w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9, N162, N163, N164, N165, N166, N167, N168, N169, N178, 
        N179, N180, N181, N182, N183, N184, N185, N194, N195, 
        N196, N197, N198, N199, N200, N201, N210, N211, N212, 
        N213, N214, N215, N216, N217, N34, N35, N36, N37, 
        N38, N388, N39, N390, N40, N404, N405, N406, N407, 
        N408, N41, N418, N419, N420, N421, N423, N425, N435, 
        N436, N437, N438, N439, N440, N441, N450, N451, N452, 
        N453, N454, N455, N456, N466, N467, N468, N469, N473, 
        N482, N483, N484, N485, N489, N498, N499, N50, N500, 
        N501, N502, N503, N504, N505, N51, N52, N53, N54, 
        N55, N56, N57, N66, N67, N68, N69, N70, N71, 
        N72, N73, N82, N83, N84, N85, N86, N87, N88, 
        N89, n1214, n1217, n1218, u0_n113, u0_n115, u0_n116, u0_n118, u0_n119, 
        u0_n121, u0_n122, u0_n124, u0_n128, u0_n130, u0_n168, u0_n174, u0_n194, u0_n196, 
        u0_n198, u0_n200, u0_n204, u0_n74, u0_n76, u0_n83, u0_n85 );
  input n1, n11, n1109, n1114, n1212, n1213, n1215, n1216, n1219, 
        n1220, n1221, n129, n13, n131, n133, n135, n137, n139, 
        n141, n143, n145, n147, n149, n15, n151, n153, n155, 
        n157, n159, n161, n163, n165, n167, n169, n17, n171, 
        n173, n175, n177, n179, n181, n183, n185, n187, n189, 
        n19, n191, n21, n23, n25, n27, n29, n3, n31, 
        n33, n35, n37, n39, n41, n43, n45, n47, n49, 
        n5, n51, n53, n55, n57, n59, n61, n63, n7, 
        n9, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, 
        sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa11_sr_0, 
        sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa13_sr_0, sa13_sr_1, 
        sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, 
        sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, 
        sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, 
        sa31_sr_5, sa31_sr_6, sa31_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, 
        sa33_sr_6, sa33_sr_7, u0_n13, u0_n250, u0_n254, u0_n258, u0_n264, u0_n33, u0_n35, 
        u0_n37, u0_n39, u0_n43, u0_n7, w1_0, w1_1, w1_10, w1_11, w1_12, 
        w1_13, w1_14, w1_15, w1_16, w1_17, w1_18, w1_19, w1_2, w1_20, 
        w1_21, w1_22, w1_23, w1_24, w1_25, w1_26, w1_27, w1_28, w1_29, 
        w1_3, w1_30, w1_31, w1_4, w1_5, w1_6, w1_7, w1_8, w1_9, 
        w2_10, w2_12, w2_13, w2_14, w2_15, w2_25, w2_28, w3_0, w3_1, 
        w3_10, w3_11, w3_16, w3_17, w3_18, w3_19, w3_2, w3_20, w3_21, 
        w3_22, w3_23, w3_24, w3_25, w3_26, w3_27, w3_28, w3_29, w3_3, 
        w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, w3_9;
  output N162, N163, N164, N165, N166, N167, N168, N169, N178, 
        N179, N180, N181, N182, N183, N184, N185, N194, N195, 
        N196, N197, N198, N199, N200, N201, N210, N211, N212, 
        N213, N214, N215, N216, N217, N34, N35, N36, N37, 
        N38, N388, N39, N390, N40, N404, N405, N406, N407, 
        N408, N41, N418, N419, N420, N421, N423, N425, N435, 
        N436, N437, N438, N439, N440, N441, N450, N451, N452, 
        N453, N454, N455, N456, N466, N467, N468, N469, N473, 
        N482, N483, N484, N485, N489, N498, N499, N50, N500, 
        N501, N502, N503, N504, N505, N51, N52, N53, N54, 
        N55, N56, N57, N66, N67, N68, N69, N70, N71, 
        N72, N73, N82, N83, N84, N85, N86, N87, N88, 
        N89, n1214, n1217, n1218, u0_n113, u0_n115, u0_n116, u0_n118, u0_n119, 
        u0_n121, u0_n122, u0_n124, u0_n128, u0_n130, u0_n168, u0_n174, u0_n194, u0_n196, 
        u0_n198, u0_n200, u0_n204, u0_n74, u0_n76, u0_n83, u0_n85;
  wire n1115, n1116, n1119, n1120, n1121, n1122, n1123, n1124, n1125, 
       n1129, n1134, n1137, n1140, n1141, n1142, n1143, n1146, n1147, 
       n1152, n1157, n1159, n1162, n1163, n1165, n1167, n1170, n1171, 
       n1174, n1175, n1176, n1177, n1180, n1182, n1184, n1185, n1187, 
       n1189, n1190, n1193, n1195, n1197, n1198, n1199, n1200, n1201, 
       n1202, n1205, n1207, n285, n286, n288, n289, n290, n291, 
       n292, n294, n295, n296, n297, n298, n300, n301, n302, 
       n303, n304, n305, n306, n307, n308, n309, n310, n311, 
       n312, n314, n315, n316, n317, n318, n319, n321, n322, 
       n323, n324, n325, n327, n328, n329, n330, n331, n332, 
       n334, n335, n336, n337, n338, n339, n341, n342, n343, 
       n345, n347, n348, n349, n350, n351, n352, n353, n354, 
       n355, n356, n357, n358, n359, n360, n361, n362, n363, 
       n365, n366, n367, n368, n369, n370, n372, n373, n374, 
       n375, n376, n378, n379, n380, n381, n382, n384, n385, 
       n386, n387, n388, n390, n391, n392, n394, n395, n396, 
       n398, n399, n400, n401, n402, n403, n404, n405, n407, 
       n408, n409, n410, n412, n413, n414, n416, n417, n418, 
       n419, n421, n422, n423, n424, n425, n426, n427, n428, 
       n429, n431, n432, n433, n434, n436, n437, n438, n439, 
       n440, n441, n442, n443, n444, n445, n446, n448, n449, 
       n450, n451, n452, n453, n454, n455, n456, n457, n459, 
       n460, n461, n462, n464, n639, n640, n642, n643, n644, 
       n645, n646, n647, n649, n650, n651, n652, n653, n655, 
       n656, n657, n658, n659, n660, n661, n662, n663, n664, 
       n665, n666, n667, n669, n670, n671, n672, n673, n674, 
       n676, n677, n678, n679, n680, n682, n683, n684, n685, 
       n686, n687, n689, n690, n691, n692, n693, n694, n696, 
       n697, n698, n700, n702, n703, n704, n705, n706, n707, 
       n708, n709, n710, n711, n712, n713, n714, n715, n716, 
       n718, n719, n720, n721, n722, n724, n725, n726, n728, 
       n729, n730, n731, n732, n734, n735, n736, n738, n739, 
       n740, n742, n743, n744, n745, n746, n747, n748, n749, 
       n750, n751, n752, n753, n755, n756, n757, n758, n760, 
       n761, n762, n764, n765, n766, n767, n769, n770, n771, 
       n772, n773, n774, n775, n776, n777, n778, n779, n780, 
       n781, n782, n783, n784, n785, n786, n787, n788, n789, 
       n790, n791, n792, n793, n794, n796, n797, n798, n799, 
       n800, n801, n802, n803, n804, n806, n807, n808, n809, 
       n810, n812, w3_12, w3_13, w3_14,  w3_15;
  XOR2_X1 U1001 (.Z( n728 ) , .B( n729 ) , .A( sa11_sr_0 ) );
  XOR2_X1 U1002 (.Z( n729 ) , .B( sa21_sr_0 ) , .A( w1_17 ) );
  XNOR2_X1 U1004 (.B( n683 ) , .ZN( n730 ) , .A( sa01_sr_1 ) );
  XOR2_X1 U1005 (.A( n163 ) , .Z( n725 ) , .B( w1_17 ) );
  OAI22_X1 U1007 (.ZN( N194 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n731 ) , .B1( n732 ) );
  XOR2_X1 U1009 (.A( n690 ) , .B( n713 ) , .Z( n734 ) );
  XOR2_X1 U1010 (.Z( n713 ) , .A( sa11_sr_7 ) , .B( sa21_sr_7 ) );
  XOR2_X1 U1012 (.A( n161 ) , .Z( n731 ) , .B( w1_16 ) );
  OAI22_X1 U1014 (.ZN( N185 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n735 ) , .B1( n736 ) );
  XOR2_X1 U1016 (.A( n650 ) , .B( n665 ) , .Z( n738 ) );
  XOR2_X1 U1017 (.Z( n650 ) , .A( sa21_sr_6 ) , .B( sa31_sr_6 ) );
  XOR2_X1 U1019 (.A( n159 ) , .Z( n735 ) , .B( w1_15 ) );
  OAI22_X1 U1021 (.ZN( N184 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n739 ) , .B1( n740 ) );
  XOR2_X1 U1023 (.A( n644 ) , .B( n656 ) , .Z( n742 ) );
  XOR2_X1 U1024 (.Z( n656 ) , .A( sa21_sr_5 ) , .B( sa31_sr_5 ) );
  XOR2_X1 U1026 (.A( n157 ) , .Z( n739 ) , .B( w1_14 ) );
  OAI22_X1 U1028 (.ZN( N183 ) , .A1( n1109 ) , .B2( n1221 ) , .A2( n743 ) , .B1( n744 ) );
  XOR2_X1 U1029 (.Z( n744 ) , .A( n745 ) , .B( n746 ) );
  XOR2_X1 U1030 (.A( n651 ) , .B( n663 ) , .Z( n746 ) );
  XOR2_X1 U1031 (.Z( n663 ) , .A( sa21_sr_4 ) , .B( sa31_sr_4 ) );
  XNOR2_X1 U1032 (.ZN( n745 ) , .B( sa31_sr_5 ) , .A( w1_13 ) );
  XOR2_X1 U1033 (.A( n155 ) , .Z( n743 ) , .B( w1_13 ) );
  OAI22_X1 U1035 (.ZN( N182 ) , .A1( n1213 ) , .B2( n1221 ) , .A2( n747 ) , .B1( n748 ) );
  XOR2_X1 U1036 (.Z( n748 ) , .A( n749 ) , .B( n750 ) );
  XOR2_X1 U1037 (.A( n657 ) , .B( n670 ) , .Z( n750 ) );
  XOR2_X1 U1038 (.Z( n670 ) , .A( sa21_sr_3 ) , .B( sa31_sr_3 ) );
  XOR2_X1 U1039 (.B( n643 ) , .Z( n749 ) , .A( n751 ) );
  XNOR2_X1 U1040 (.ZN( n751 ) , .B( sa31_sr_4 ) , .A( w1_12 ) );
  XOR2_X1 U1041 (.A( n153 ) , .Z( n747 ) , .B( w1_12 ) );
  OAI22_X1 U1043 (.ZN( N181 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n752 ) , .B1( n753 ) );
  XOR2_X1 U1045 (.A( n662 ) , .B( n677 ) , .Z( n755 ) );
  XOR2_X1 U1046 (.Z( n677 ) , .A( sa21_sr_2 ) , .B( sa31_sr_2 ) );
  XNOR2_X1 U1048 (.ZN( n756 ) , .B( sa31_sr_3 ) , .A( w1_11 ) );
  XOR2_X1 U1049 (.A( n151 ) , .Z( n752 ) , .B( w1_11 ) );
  OAI22_X1 U1051 (.ZN( N180 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n757 ) , .B1( n758 ) );
  XOR2_X1 U1053 (.A( n671 ) , .B( n683 ) , .Z( n760 ) );
  XOR2_X1 U1054 (.Z( n683 ) , .A( sa21_sr_1 ) , .B( sa31_sr_1 ) );
  XOR2_X1 U1056 (.A( n149 ) , .Z( n757 ) , .B( w1_10 ) );
  OAI22_X1 U1058 (.ZN( N179 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n761 ) , .B1( n762 ) );
  XOR2_X1 U1060 (.A( n678 ) , .B( n690 ) , .Z( n764 ) );
  XOR2_X1 U1061 (.Z( n690 ) , .A( sa21_sr_0 ) , .B( sa31_sr_0 ) );
  XNOR2_X1 U1063 (.ZN( n765 ) , .B( sa31_sr_1 ) , .A( w1_9 ) );
  XOR2_X1 U1064 (.A( n147 ) , .Z( n761 ) , .B( w1_9 ) );
  OAI22_X1 U1066 (.ZN( N178 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n766 ) , .B1( n767 ) );
  XOR2_X1 U1068 (.A( n643 ) , .B( n684 ) , .Z( n769 ) );
  XOR2_X1 U1069 (.Z( n643 ) , .A( sa21_sr_7 ) , .B( sa31_sr_7 ) );
  XOR2_X1 U1071 (.A( n145 ) , .Z( n766 ) , .B( w1_8 ) );
  OAI22_X1 U1073 (.ZN( N169 ) , .A1( n1109 ) , .B2( n1217 ) , .A2( n770 ) , .B1( n771 ) );
  XOR2_X1 U1074 (.Z( n771 ) , .A( n772 ) , .B( n773 ) );
  XOR2_X1 U1075 (.B( n665 ) , .Z( n773 ) , .A( sa01_sr_6 ) );
  XOR2_X1 U1076 (.Z( n665 ) , .A( sa01_sr_7 ) , .B( sa11_sr_7 ) );
  XNOR2_X1 U1077 (.ZN( n772 ) , .B( n774 ) , .A( sa21_sr_7 ) );
  XOR2_X1 U1078 (.Z( n774 ) , .B( sa31_sr_6 ) , .A( w1_7 ) );
  XOR2_X1 U1079 (.A( n143 ) , .Z( n770 ) , .B( w1_7 ) );
  OAI22_X1 U1081 (.ZN( N168 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n775 ) , .B1( n776 ) );
  XOR2_X1 U1082 (.Z( n776 ) , .A( n777 ) , .B( n778 ) );
  XOR2_X1 U1083 (.Z( n778 ) , .B( n779 ) , .A( sa21_sr_6 ) );
  XOR2_X1 U1084 (.Z( n779 ) , .B( sa31_sr_5 ) , .A( w1_6 ) );
  XNOR2_X1 U1085 (.B( n644 ) , .ZN( n777 ) , .A( sa01_sr_5 ) );
  XOR2_X1 U1086 (.Z( n644 ) , .A( sa01_sr_6 ) , .B( sa11_sr_6 ) );
  XOR2_X1 U1087 (.A( n141 ) , .Z( n775 ) , .B( w1_6 ) );
  OAI22_X1 U1089 (.ZN( N167 ) , .A1( n1212 ) , .B2( n1217 ) , .A2( n780 ) , .B1( n781 ) );
  XOR2_X1 U1090 (.Z( n781 ) , .A( n782 ) , .B( n783 ) );
  XOR2_X1 U1091 (.Z( n783 ) , .B( n784 ) , .A( sa21_sr_5 ) );
  XOR2_X1 U1092 (.Z( n784 ) , .B( sa31_sr_4 ) , .A( w1_5 ) );
  XNOR2_X1 U1093 (.B( n651 ) , .ZN( n782 ) , .A( sa01_sr_4 ) );
  XOR2_X1 U1094 (.Z( n651 ) , .A( sa01_sr_5 ) , .B( sa11_sr_5 ) );
  XOR2_X1 U1095 (.A( n139 ) , .Z( n780 ) , .B( w1_5 ) );
  OAI22_X1 U1097 (.ZN( N166 ) , .A1( n1213 ) , .B2( n1220 ) , .A2( n785 ) , .B1( n786 ) );
  XOR2_X1 U1098 (.Z( n786 ) , .A( n787 ) , .B( n788 ) );
  XOR2_X1 U1099 (.Z( n788 ) , .B( n789 ) , .A( sa21_sr_4 ) );
  XOR2_X1 U1100 (.Z( n789 ) , .B( sa31_sr_3 ) , .A( w1_4 ) );
  XOR2_X1 U1101 (.Z( n787 ) , .A( n790 ) , .B( n791 ) );
  XNOR2_X1 U1102 (.B( n657 ) , .ZN( n790 ) , .A( sa01_sr_3 ) );
  XOR2_X1 U1103 (.Z( n657 ) , .A( sa01_sr_4 ) , .B( sa11_sr_4 ) );
  XOR2_X1 U1104 (.A( n137 ) , .Z( n785 ) , .B( w1_4 ) );
  OAI22_X1 U1106 (.ZN( N165 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n792 ) , .B1( n793 ) );
  XOR2_X1 U1109 (.Z( n796 ) , .B( sa31_sr_2 ) , .A( w1_3 ) );
  XOR2_X1 U1110 (.B( n791 ) , .Z( n794 ) , .A( n797 ) );
  XNOR2_X1 U1111 (.B( n662 ) , .ZN( n797 ) , .A( sa01_sr_2 ) );
  XOR2_X1 U1112 (.Z( n662 ) , .A( sa01_sr_3 ) , .B( sa11_sr_3 ) );
  XOR2_X1 U1113 (.A( n135 ) , .Z( n792 ) , .B( w1_3 ) );
  OAI22_X1 U1115 (.ZN( N164 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n798 ) , .B1( n799 ) );
  XOR2_X1 U1116 (.Z( n799 ) , .A( n800 ) , .B( n801 ) );
  XOR2_X1 U1117 (.Z( n801 ) , .B( n802 ) , .A( sa21_sr_2 ) );
  XOR2_X1 U1118 (.Z( n802 ) , .B( sa31_sr_1 ) , .A( w1_2 ) );
  XNOR2_X1 U1119 (.B( n671 ) , .ZN( n800 ) , .A( sa01_sr_1 ) );
  XOR2_X1 U1120 (.Z( n671 ) , .A( sa01_sr_2 ) , .B( sa11_sr_2 ) );
  XOR2_X1 U1121 (.A( n133 ) , .Z( n798 ) , .B( w1_2 ) );
  OAI22_X1 U1123 (.ZN( N163 ) , .A1( n1215 ) , .B2( n1220 ) , .A2( n803 ) , .B1( n804 ) );
  XOR2_X1 U1125 (.Z( n806 ) , .B( n807 ) , .A( sa21_sr_1 ) );
  XOR2_X1 U1126 (.Z( n807 ) , .B( sa31_sr_0 ) , .A( w1_1 ) );
  XNOR2_X1 U1128 (.B( n678 ) , .ZN( n808 ) , .A( sa01_sr_0 ) );
  XOR2_X1 U1129 (.Z( n678 ) , .A( sa01_sr_1 ) , .B( sa11_sr_1 ) );
  XOR2_X1 U1130 (.A( n131 ) , .Z( n803 ) , .B( w1_1 ) );
  OAI22_X1 U1132 (.ZN( N162 ) , .A1( n1215 ) , .B2( n1217 ) , .A2( n809 ) , .B1( n810 ) );
  XOR2_X1 U1134 (.A( n684 ) , .B( n791 ) , .Z( n812 ) );
  XOR2_X1 U1135 (.Z( n791 ) , .A( sa01_sr_7 ) , .B( sa31_sr_7 ) );
  XOR2_X1 U1136 (.Z( n684 ) , .A( sa01_sr_0 ) , .B( sa11_sr_0 ) );
  XOR2_X1 U1138 (.A( n129 ) , .Z( n809 ) , .B( w1_0 ) );
  XOR2_X1 U1370 (.A( n1115 ) , .Z( n382 ) , .B( n384 ) );
  XOR2_X1 U1371 (.Z( n1115 ) , .B( n386 ) , .A( w3_16 ) );
  XNOR2_X1 U1372 (.B( n1116 ) , .ZN( n338 ) , .A( sa13_sr_6 ) );
  XOR2_X1 U1373 (.Z( n1116 ) , .B( sa23_sr_6 ) , .A( w3_23 ) );
  XNOR2_X1 U1381 (.B( n650 ) , .ZN( n698 ) , .A( sa01_sr_6 ) );
  XNOR2_X1 U1382 (.B( n295 ) , .ZN( n343 ) , .A( sa03_sr_6 ) );
  INV_X1 U1384 (.A( n1114 ) , .ZN( n1214 ) );
  BUF_X1 U1385 (.Z( n1217 ) , .A( n1221 ) );
  BUF_X1 U1386 (.Z( n1218 ) , .A( n1221 ) );
  XNOR2_X1 U1387 (.A( n1119 ) , .ZN( n405 ) , .B( n407 ) );
  XNOR2_X1 U1388 (.ZN( n1119 ) , .B( n289 ) , .A( n408 ) );
  XNOR2_X1 U1389 (.A( n1120 ) , .ZN( n312 ) , .B( n314 ) );
  XNOR2_X1 U1390 (.ZN( n1120 ) , .B( n307 ) , .A( n317 ) );
  XNOR2_X1 U1391 (.A( n1121 ) , .ZN( n392 ) , .B( n394 ) );
  XOR2_X1 U1392 (.Z( n1121 ) , .B( sa33_sr_6 ) , .A( w3_14 ) );
  XNOR2_X1 U1393 (.B( n1122 ) , .ZN( n428 ) , .A( n429 ) );
  XNOR2_X1 U1394 (.ZN( n1122 ) , .B( n431 ) , .A( sa23_sr_6 ) );
  XNOR2_X1 U1395 (.A( n1123 ) , .ZN( n388 ) , .B( n390 ) );
  XOR2_X1 U1396 (.Z( n1123 ) , .B( sa33_sr_7 ) , .A( w3_15 ) );
  XNOR2_X1 U1397 (.A( n1124 ) , .ZN( n396 ) , .B( n398 ) );
  XOR2_X1 U1398 (.Z( n1124 ) , .B( sa33_sr_5 ) , .A( w3_13 ) );
  XNOR2_X1 U1401 (.A( n1125 ) , .ZN( n753 ) , .B( n755 ) );
  XNOR2_X1 U1402 (.ZN( n1125 ) , .B( n643 ) , .A( n756 ) );
  XNOR2_X1 U1409 (.A( n1129 ) , .ZN( n667 ) , .B( n669 ) );
  XNOR2_X1 U1410 (.ZN( n1129 ) , .B( n665 ) , .A( n672 ) );
  XNOR2_X1 U1419 (.B( n1134 ) , .ZN( n433 ) , .A( n434 ) );
  XNOR2_X1 U1420 (.ZN( n1134 ) , .B( n436 ) , .A( sa23_sr_5 ) );
  XNOR2_X1 U1425 (.A( n1137 ) , .ZN( n325 ) , .B( n327 ) );
  XNOR2_X1 U1426 (.ZN( n1137 ) , .B( n307 ) , .A( n330 ) );
  XNOR2_X1 U1431 (.B( n1140 ) , .ZN( n445 ) , .A( n446 ) );
  XNOR2_X1 U1432 (.ZN( n1140 ) , .B( n448 ) , .A( sa23_sr_3 ) );
  XNOR2_X1 U1433 (.B( n1141 ) , .ZN( n362 ) , .A( n363 ) );
  XNOR2_X1 U1434 (.ZN( n1141 ) , .B( n365 ) , .A( sa13_sr_2 ) );
  XNOR2_X1 U1435 (.B( n1142 ) , .ZN( n369 ) , .A( n370 ) );
  XNOR2_X1 U1436 (.ZN( n1142 ) , .B( n372 ) , .A( sa13_sr_1 ) );
  XNOR2_X1 U1437 (.B( n1143 ) , .ZN( n715 ) , .A( n716 ) );
  XNOR2_X1 U1438 (.ZN( n1143 ) , .B( n718 ) , .A( sa11_sr_2 ) );
  XNOR2_X1 U1443 (.A( n1146 ) , .ZN( n640 ) , .B( n642 ) );
  XNOR2_X1 U1444 (.ZN( n1146 ) , .B( n645 ) , .A( w1_31 ) );
  XNOR2_X1 U1445 (.A( n1147 ) , .ZN( n687 ) , .B( n689 ) );
  XOR2_X1 U1446 (.Z( n1147 ) , .B( sa11_sr_0 ) , .A( w1_24 ) );
  XNOR2_X1 U1455 (.A( n1152 ) , .ZN( n736 ) , .B( n738 ) );
  XOR2_X1 U1456 (.Z( n1152 ) , .B( sa31_sr_7 ) , .A( w1_15 ) );
  XNOR2_X1 U1465 (.A( n1157 ) , .ZN( n647 ) , .B( n649 ) );
  XOR2_X1 U1466 (.Z( n1157 ) , .B( sa11_sr_6 ) , .A( w1_30 ) );
  XNOR2_X1 U1469 (.A( n1159 ) , .ZN( n762 ) , .B( n764 ) );
  XNOR2_X1 U1470 (.ZN( n1159 ) , .B( n643 ) , .A( n765 ) );
  XNOR2_X1 U1475 (.B( n1162 ) , .ZN( n697 ) , .A( n698 ) );
  XNOR2_X1 U1476 (.ZN( n1162 ) , .B( n700 ) , .A( sa11_sr_5 ) );
  XNOR2_X1 U1477 (.A( n1163 ) , .ZN( n740 ) , .B( n742 ) );
  XOR2_X1 U1478 (.Z( n1163 ) , .B( sa31_sr_6 ) , .A( w1_14 ) );
  XNOR2_X1 U1481 (.A( n1165 ) , .ZN( n414 ) , .B( n416 ) );
  XNOR2_X1 U1482 (.ZN( n1165 ) , .B( n289 ) , .A( n417 ) );
  XNOR2_X1 U1485 (.B( n1167 ) , .ZN( n793 ) , .A( n794 ) );
  XNOR2_X1 U1486 (.ZN( n1167 ) , .B( n796 ) , .A( sa21_sr_3 ) );
  XNOR2_X1 U1491 (.A( n1170 ) , .ZN( n767 ) , .B( n769 ) );
  XOR2_X1 U1492 (.Z( n1170 ) , .B( sa31_sr_0 ) , .A( w1_8 ) );
  XNOR2_X1 U1493 (.A( n1171 ) , .ZN( n732 ) , .B( n734 ) );
  XOR2_X1 U1494 (.Z( n1171 ) , .B( sa01_sr_0 ) , .A( w1_16 ) );
  XNOR2_X1 U1499 (.A( n1174 ) , .ZN( n653 ) , .B( n655 ) );
  XOR2_X1 U1500 (.Z( n1174 ) , .B( sa11_sr_5 ) , .A( w1_29 ) );
  XNOR2_X1 U1501 (.B( n1175 ) , .ZN( n456 ) , .A( n457 ) );
  XNOR2_X1 U1502 (.ZN( n1175 ) , .B( n459 ) , .A( sa23_sr_1 ) );
  XNOR2_X1 U1503 (.B( n1176 ) , .ZN( n721 ) , .A( n722 ) );
  XNOR2_X1 U1504 (.ZN( n1176 ) , .B( n724 ) , .A( sa11_sr_1 ) );
  XNOR2_X1 U1505 (.A( n1177 ) , .ZN( n680 ) , .B( n682 ) );
  XNOR2_X1 U1506 (.ZN( n1177 ) , .B( n665 ) , .A( n685 ) );
  XNOR2_X1 U1511 (.B( n1180 ) , .ZN( n375 ) , .A( n376 ) );
  XNOR2_X1 U1512 (.ZN( n1180 ) , .B( n378 ) , .A( sa13_sr_0 ) );
  XNOR2_X1 U1515 (.B( n1182 ) , .ZN( n342 ) , .A( n343 ) );
  XNOR2_X1 U1516 (.ZN( n1182 ) , .B( n345 ) , .A( sa13_sr_5 ) );
  XNOR2_X1 U1519 (.A( n1184 ) , .ZN( n810 ) , .B( n812 ) );
  XOR2_X1 U1520 (.Z( n1184 ) , .B( sa21_sr_0 ) , .A( w1_0 ) );
  XNOR2_X1 U1521 (.A( n1185 ) , .ZN( n726 ) , .B( n728 ) );
  XNOR2_X1 U1522 (.ZN( n1185 ) , .B( n713 ) , .A( n730 ) );
  XNOR2_X1 U1525 (.A( n1187 ) , .ZN( n804 ) , .B( n806 ) );
  XNOR2_X1 U1526 (.ZN( n1187 ) , .B( n791 ) , .A( n808 ) );
  XOR2_X1 U1529 (.B( n1189 ) , .Z( n693 ) , .A( sa11_sr_6 ) );
  XNOR2_X1 U1530 (.ZN( n1189 ) , .B( sa21_sr_6 ) , .A( w1_23 ) );
  XNOR2_X1 U1531 (.A( n1190 ) , .ZN( n419 ) , .B( n421 ) );
  XOR2_X1 U1532 (.Z( n1190 ) , .B( sa33_sr_0 ) , .A( w3_8 ) );
  XNOR2_X1 U1537 (.A( n1193 ) , .ZN( n332 ) , .B( n334 ) );
  XOR2_X1 U1538 (.Z( n1193 ) , .B( sa13_sr_0 ) , .A( w3_24 ) );
  XNOR2_X1 U1541 (.A( n1195 ) , .ZN( n286 ) , .B( n288 ) );
  XOR2_X1 U1542 (.Z( n1195 ) , .B( sa13_sr_7 ) , .A( w3_31 ) );
  XNOR2_X1 U1545 (.A( n1197 ) , .ZN( n674 ) , .B( n676 ) );
  XOR2_X1 U1546 (.Z( n1197 ) , .B( sa11_sr_2 ) , .A( w1_26 ) );
  XNOR2_X1 U1547 (.A( n1198 ) , .ZN( n758 ) , .B( n760 ) );
  XOR2_X1 U1548 (.Z( n1198 ) , .B( sa31_sr_2 ) , .A( w1_10 ) );
  XNOR2_X1 U1549 (.A( n1199 ) , .ZN( n298 ) , .B( n300 ) );
  XOR2_X1 U1550 (.Z( n1199 ) , .B( sa13_sr_5 ) , .A( w3_29 ) );
  XNOR2_X1 U1551 (.A( n1200 ) , .ZN( n319 ) , .B( n321 ) );
  XOR2_X1 U1552 (.Z( n1200 ) , .B( sa13_sr_2 ) , .A( w3_26 ) );
  XNOR2_X1 U1553 (.A( n1201 ) , .ZN( n410 ) , .B( n412 ) );
  XOR2_X1 U1554 (.Z( n1201 ) , .B( sa33_sr_2 ) , .A( w3_10 ) );
  XNOR2_X1 U1555 (.A( n1202 ) , .ZN( n462 ) , .B( n464 ) );
  XOR2_X1 U1556 (.Z( n1202 ) , .B( sa23_sr_0 ) , .A( w3_0 ) );
  XNOR2_X1 U1561 (.A( n1205 ) , .ZN( n292 ) , .B( n294 ) );
  XOR2_X1 U1562 (.Z( n1205 ) , .B( sa13_sr_6 ) , .A( w3_30 ) );
  XNOR2_X1 U1566 (.ZN( N423 ) , .B( n1207 ) , .A( w1_18 ) );
  INV_X1 U1568 (.ZN( n1207 ) , .A( sa11_sr_2 ) );
  OAI22_X1 U290 (.ZN( N89 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n285 ) , .B1( n286 ) );
  XOR2_X1 U292 (.Z( n288 ) , .A( n289 ) , .B( n290 ) );
  XOR2_X1 U294 (.Z( n285 ) , .A( n63 ) , .B( w3_31 ) );
  OAI22_X1 U296 (.ZN( N88 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n291 ) , .B1( n292 ) );
  XOR2_X1 U298 (.Z( n294 ) , .A( n295 ) , .B( n296 ) );
  XOR2_X1 U300 (.Z( n291 ) , .A( n61 ) , .B( w3_30 ) );
  OAI22_X1 U302 (.ZN( N87 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n297 ) , .B1( n298 ) );
  XOR2_X1 U304 (.Z( n300 ) , .A( n301 ) , .B( n302 ) );
  XOR2_X1 U306 (.Z( n297 ) , .A( n59 ) , .B( w3_29 ) );
  OAI22_X1 U308 (.ZN( N86 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n303 ) , .B1( n304 ) );
  XOR2_X1 U309 (.Z( n304 ) , .A( n305 ) , .B( n306 ) );
  XOR2_X1 U310 (.Z( n306 ) , .A( n307 ) , .B( n308 ) );
  XOR2_X1 U311 (.Z( n305 ) , .A( n309 ) , .B( n310 ) );
  XNOR2_X1 U312 (.ZN( n309 ) , .B( sa13_sr_4 ) , .A( w3_28 ) );
  XOR2_X1 U313 (.Z( n303 ) , .A( n57 ) , .B( w3_28 ) );
  OAI22_X1 U315 (.ZN( N85 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n311 ) , .B1( n312 ) );
  XOR2_X1 U317 (.Z( n314 ) , .A( n315 ) , .B( n316 ) );
  XNOR2_X1 U319 (.ZN( n317 ) , .B( sa13_sr_3 ) , .A( w3_27 ) );
  XOR2_X1 U320 (.Z( n311 ) , .A( n55 ) , .B( w3_27 ) );
  OAI22_X1 U322 (.ZN( N84 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n318 ) , .B1( n319 ) );
  XOR2_X1 U324 (.Z( n321 ) , .A( n322 ) , .B( n323 ) );
  XOR2_X1 U326 (.Z( n318 ) , .A( n53 ) , .B( w3_26 ) );
  OAI22_X1 U328 (.ZN( N83 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n324 ) , .B1( n325 ) );
  XOR2_X1 U330 (.Z( n327 ) , .A( n328 ) , .B( n329 ) );
  XNOR2_X1 U332 (.ZN( n330 ) , .B( sa13_sr_1 ) , .A( w3_25 ) );
  XOR2_X1 U333 (.Z( n324 ) , .A( n51 ) , .B( w3_25 ) );
  OAI22_X1 U335 (.ZN( N82 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n331 ) , .B1( n332 ) );
  XOR2_X1 U337 (.A( n307 ) , .Z( n334 ) , .B( n335 ) );
  XOR2_X1 U339 (.Z( n331 ) , .A( n49 ) , .B( w3_24 ) );
  OAI22_X1 U341 (.ZN( N73 ) , .A1( n1213 ) , .B2( n1219 ) , .A2( n336 ) , .B1( n337 ) );
  XOR2_X1 U342 (.Z( n337 ) , .A( n338 ) , .B( n339 ) );
  XOR2_X1 U343 (.B( n289 ) , .Z( n339 ) , .A( sa03_sr_7 ) );
  XOR2_X1 U346 (.Z( n336 ) , .A( n47 ) , .B( w3_23 ) );
  OAI22_X1 U348 (.ZN( N72 ) , .A1( n1212 ) , .B2( n1217 ) , .A2( n341 ) , .B1( n342 ) );
  XOR2_X1 U351 (.Z( n345 ) , .B( sa23_sr_5 ) , .A( w3_22 ) );
  XOR2_X1 U354 (.Z( n341 ) , .A( n45 ) , .B( w3_22 ) );
  OAI22_X1 U356 (.ZN( N71 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n347 ) , .B1( n348 ) );
  XOR2_X1 U357 (.Z( n348 ) , .A( n349 ) , .B( n350 ) );
  XOR2_X1 U358 (.Z( n350 ) , .B( n351 ) , .A( sa13_sr_4 ) );
  XOR2_X1 U359 (.Z( n351 ) , .B( sa23_sr_4 ) , .A( w3_21 ) );
  XOR2_X1 U360 (.B( n301 ) , .Z( n349 ) , .A( n352 ) );
  XOR2_X1 U361 (.Z( n347 ) , .A( n43 ) , .B( w3_21 ) );
  OAI22_X1 U363 (.ZN( N70 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n353 ) , .B1( n354 ) );
  XOR2_X1 U364 (.Z( n354 ) , .A( n355 ) , .B( n356 ) );
  XOR2_X1 U365 (.Z( n356 ) , .B( n357 ) , .A( sa13_sr_3 ) );
  XOR2_X1 U366 (.Z( n357 ) , .B( sa23_sr_3 ) , .A( w3_20 ) );
  XOR2_X1 U367 (.Z( n355 ) , .A( n358 ) , .B( n359 ) );
  XOR2_X1 U368 (.B( n310 ) , .Z( n358 ) , .A( n360 ) );
  XOR2_X1 U369 (.Z( n353 ) , .A( n41 ) , .B( w3_20 ) );
  OAI22_X1 U371 (.ZN( N69 ) , .B2( n1114 ) , .A1( n1212 ) , .A2( n361 ) , .B1( n362 ) );
  XOR2_X1 U374 (.Z( n365 ) , .B( sa23_sr_2 ) , .A( w3_19 ) );
  XOR2_X1 U375 (.B( n359 ) , .Z( n363 ) , .A( n366 ) );
  XOR2_X1 U376 (.B( n315 ) , .Z( n366 ) , .A( n367 ) );
  XOR2_X1 U377 (.Z( n361 ) , .A( n39 ) , .B( w3_19 ) );
  OAI22_X1 U379 (.ZN( N68 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n368 ) , .B1( n369 ) );
  XOR2_X1 U382 (.Z( n372 ) , .B( sa23_sr_1 ) , .A( w3_18 ) );
  XOR2_X1 U383 (.B( n322 ) , .Z( n370 ) , .A( n373 ) );
  XOR2_X1 U384 (.Z( n368 ) , .A( n37 ) , .B( w3_18 ) );
  OAI22_X1 U386 (.ZN( N67 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n374 ) , .B1( n375 ) );
  XOR2_X1 U389 (.Z( n378 ) , .B( sa23_sr_0 ) , .A( w3_17 ) );
  XOR2_X1 U390 (.B( n359 ) , .Z( n376 ) , .A( n379 ) );
  XOR2_X1 U391 (.B( n328 ) , .Z( n379 ) , .A( n380 ) );
  XOR2_X1 U392 (.A( n35 ) , .Z( n374 ) , .B( w3_17 ) );
  OAI22_X1 U394 (.ZN( N66 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n381 ) , .B1( n382 ) );
  XOR2_X1 U396 (.A( n335 ) , .B( n359 ) , .Z( n384 ) );
  XNOR2_X1 U397 (.ZN( n359 ) , .B( n385 ) , .A( sa13_sr_7 ) );
  XOR2_X1 U399 (.A( n33 ) , .Z( n381 ) , .B( w3_16 ) );
  OAI22_X1 U401 (.ZN( N57 ) , .A1( n1212 ) , .B2( n1221 ) , .A2( n387 ) , .B1( n388 ) );
  XOR2_X1 U403 (.A( n295 ) , .B( n307 ) , .Z( n390 ) );
  XOR2_X1 U404 (.Z( n295 ) , .A( sa23_sr_6 ) , .B( sa33_sr_6 ) );
  XOR2_X1 U406 (.A( n31 ) , .Z( n387 ) , .B( w3_15 ) );
  OAI22_X1 U408 (.ZN( N56 ) , .B2( n1114 ) , .A1( n1213 ) , .A2( n391 ) , .B1( n392 ) );
  XOR2_X1 U410 (.A( n290 ) , .B( n301 ) , .Z( n394 ) );
  XOR2_X1 U411 (.Z( n301 ) , .A( sa23_sr_5 ) , .B( sa33_sr_5 ) );
  XOR2_X1 U413 (.A( n29 ) , .Z( n391 ) , .B( w3_14 ) );
  OAI22_X1 U415 (.ZN( N55 ) , .A1( n1216 ) , .B2( n1221 ) , .A2( n395 ) , .B1( n396 ) );
  XOR2_X1 U417 (.A( n296 ) , .B( n310 ) , .Z( n398 ) );
  XOR2_X1 U418 (.Z( n310 ) , .A( sa23_sr_4 ) , .B( sa33_sr_4 ) );
  XOR2_X1 U420 (.A( n27 ) , .Z( n395 ) , .B( w3_13 ) );
  OAI22_X1 U422 (.ZN( N54 ) , .A1( n1216 ) , .B2( n1220 ) , .A2( n399 ) , .B1( n400 ) );
  XOR2_X1 U423 (.Z( n400 ) , .A( n401 ) , .B( n402 ) );
  XOR2_X1 U424 (.A( n302 ) , .B( n315 ) , .Z( n402 ) );
  XOR2_X1 U425 (.Z( n315 ) , .A( sa23_sr_3 ) , .B( sa33_sr_3 ) );
  XOR2_X1 U426 (.B( n289 ) , .Z( n401 ) , .A( n403 ) );
  XNOR2_X1 U427 (.ZN( n403 ) , .B( sa33_sr_4 ) , .A( w3_12 ) );
  XOR2_X1 U428 (.A( n25 ) , .Z( n399 ) , .B( w3_12 ) );
  OAI22_X1 U430 (.ZN( N53 ) , .A1( n1216 ) , .B2( n1220 ) , .A2( n404 ) , .B1( n405 ) );
  XOR2_X1 U432 (.A( n308 ) , .B( n322 ) , .Z( n407 ) );
  XOR2_X1 U433 (.Z( n322 ) , .A( sa23_sr_2 ) , .B( sa33_sr_2 ) );
  XNOR2_X1 U435 (.ZN( n408 ) , .B( sa33_sr_3 ) , .A( w3_11 ) );
  XOR2_X1 U436 (.A( n23 ) , .Z( n404 ) , .B( w3_11 ) );
  OAI22_X1 U438 (.ZN( N52 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n409 ) , .B1( n410 ) );
  XOR2_X1 U440 (.A( n316 ) , .B( n328 ) , .Z( n412 ) );
  XOR2_X1 U441 (.Z( n328 ) , .A( sa23_sr_1 ) , .B( sa33_sr_1 ) );
  XOR2_X1 U443 (.A( n21 ) , .Z( n409 ) , .B( w3_10 ) );
  OAI22_X1 U445 (.ZN( N51 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n413 ) , .B1( n414 ) );
  XOR2_X1 U447 (.A( n323 ) , .B( n335 ) , .Z( n416 ) );
  XOR2_X1 U448 (.Z( n335 ) , .A( sa23_sr_0 ) , .B( sa33_sr_0 ) );
  XNOR2_X1 U450 (.ZN( n417 ) , .B( sa33_sr_1 ) , .A( w3_9 ) );
  XOR2_X1 U451 (.A( n19 ) , .Z( n413 ) , .B( w3_9 ) );
  XOR2_X1 U453 (.Z( N505 ) , .B( sa33_sr_0 ) , .A( w3_0 ) );
  XOR2_X1 U454 (.Z( N504 ) , .B( sa33_sr_1 ) , .A( w3_1 ) );
  XOR2_X1 U455 (.Z( N503 ) , .B( sa33_sr_2 ) , .A( w3_2 ) );
  XOR2_X1 U456 (.Z( N502 ) , .B( sa33_sr_3 ) , .A( w3_3 ) );
  XOR2_X1 U457 (.Z( N501 ) , .B( sa33_sr_4 ) , .A( w3_4 ) );
  XOR2_X1 U458 (.Z( N500 ) , .B( sa33_sr_5 ) , .A( w3_5 ) );
  OAI22_X1 U459 (.ZN( N50 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n418 ) , .B1( n419 ) );
  XOR2_X1 U461 (.A( n289 ) , .B( n329 ) , .Z( n421 ) );
  XOR2_X1 U462 (.Z( n289 ) , .A( sa23_sr_7 ) , .B( sa33_sr_7 ) );
  XOR2_X1 U464 (.A( n17 ) , .Z( n418 ) , .B( w3_8 ) );
  XOR2_X1 U466 (.Z( N499 ) , .B( sa33_sr_6 ) , .A( w3_6 ) );
  XOR2_X1 U467 (.Z( N498 ) , .B( sa33_sr_7 ) , .A( w3_7 ) );
  XOR2_X1 U476 (.Z( N489 ) , .B( sa31_sr_0 ) , .A( w1_0 ) );
  XOR2_X1 U480 (.Z( N485 ) , .B( sa31_sr_4 ) , .A( w1_4 ) );
  XOR2_X1 U481 (.Z( N484 ) , .B( sa31_sr_5 ) , .A( w1_5 ) );
  XOR2_X1 U482 (.Z( N483 ) , .B( sa31_sr_6 ) , .A( w1_6 ) );
  XOR2_X1 U483 (.Z( N482 ) , .B( sa31_sr_7 ) , .A( w1_7 ) );
  XOR2_X1 U492 (.Z( N473 ) , .B( sa23_sr_0 ) , .A( w3_8 ) );
  XOR2_X1 U496 (.Z( N469 ) , .B( sa23_sr_4 ) , .A( w3_12 ) );
  XOR2_X1 U497 (.Z( N468 ) , .B( sa23_sr_5 ) , .A( w3_13 ) );
  XOR2_X1 U498 (.Z( N467 ) , .B( sa23_sr_6 ) , .A( w3_14 ) );
  XOR2_X1 U499 (.Z( N466 ) , .B( sa23_sr_7 ) , .A( w3_15 ) );
  XOR2_X1 U509 (.Z( N456 ) , .B( sa21_sr_1 ) , .A( w1_9 ) );
  XOR2_X1 U510 (.Z( N455 ) , .B( sa21_sr_2 ) , .A( w1_10 ) );
  XOR2_X1 U511 (.Z( N454 ) , .B( sa21_sr_3 ) , .A( w1_11 ) );
  XOR2_X1 U512 (.Z( N453 ) , .B( sa21_sr_4 ) , .A( w1_12 ) );
  XOR2_X1 U513 (.Z( N452 ) , .B( sa21_sr_5 ) , .A( w1_13 ) );
  XOR2_X1 U514 (.Z( N451 ) , .B( sa21_sr_6 ) , .A( w1_14 ) );
  XOR2_X1 U515 (.Z( N450 ) , .B( sa21_sr_7 ) , .A( w1_15 ) );
  XOR2_X1 U524 (.Z( N441 ) , .B( sa13_sr_0 ) , .A( w3_16 ) );
  XOR2_X1 U525 (.Z( N440 ) , .B( sa13_sr_1 ) , .A( w3_17 ) );
  XOR2_X1 U526 (.Z( N439 ) , .B( sa13_sr_2 ) , .A( w3_18 ) );
  XOR2_X1 U527 (.Z( N438 ) , .B( sa13_sr_3 ) , .A( w3_19 ) );
  XOR2_X1 U528 (.Z( N437 ) , .B( sa13_sr_4 ) , .A( w3_20 ) );
  XOR2_X1 U529 (.Z( N436 ) , .B( sa13_sr_5 ) , .A( w3_21 ) );
  XOR2_X1 U530 (.Z( N435 ) , .B( sa13_sr_6 ) , .A( w3_22 ) );
  XOR2_X1 U540 (.Z( N425 ) , .B( sa11_sr_0 ) , .A( w1_16 ) );
  XOR2_X1 U544 (.Z( N421 ) , .B( sa11_sr_4 ) , .A( w1_20 ) );
  XOR2_X1 U545 (.Z( N420 ) , .B( sa11_sr_5 ) , .A( w1_21 ) );
  XOR2_X1 U546 (.Z( N419 ) , .B( sa11_sr_6 ) , .A( w1_22 ) );
  XOR2_X1 U547 (.Z( N418 ) , .B( sa11_sr_7 ) , .A( w1_23 ) );
  OAI22_X1 U556 (.ZN( N41 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n422 ) , .B1( n423 ) );
  XOR2_X1 U557 (.Z( n423 ) , .A( n424 ) , .B( n425 ) );
  XOR2_X1 U558 (.B( n307 ) , .Z( n425 ) , .A( sa03_sr_6 ) );
  XOR2_X1 U559 (.Z( n307 ) , .A( sa03_sr_7 ) , .B( sa13_sr_7 ) );
  XOR2_X1 U560 (.A( n385 ) , .Z( n424 ) , .B( n426 ) );
  XOR2_X1 U561 (.Z( n426 ) , .B( sa33_sr_6 ) , .A( w3_7 ) );
  INV_X1 U562 (.ZN( n385 ) , .A( sa23_sr_7 ) );
  XOR2_X1 U563 (.A( n15 ) , .Z( n422 ) , .B( w3_7 ) );
  XOR2_X1 U566 (.Z( N408 ) , .B( sa03_sr_1 ) , .A( w3_25 ) );
  XOR2_X1 U567 (.Z( N407 ) , .B( sa03_sr_2 ) , .A( w3_26 ) );
  XOR2_X1 U568 (.Z( N406 ) , .B( sa03_sr_3 ) , .A( w3_27 ) );
  XOR2_X1 U569 (.Z( N405 ) , .B( sa03_sr_4 ) , .A( w3_28 ) );
  XOR2_X1 U570 (.Z( N404 ) , .B( sa03_sr_5 ) , .A( w3_29 ) );
  OAI22_X1 U575 (.ZN( N40 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n427 ) , .B1( n428 ) );
  XOR2_X1 U578 (.Z( n431 ) , .B( sa33_sr_5 ) , .A( w3_6 ) );
  XOR2_X1 U579 (.B( n290 ) , .A( n352 ) , .Z( n429 ) );
  XOR2_X1 U580 (.Z( n290 ) , .A( sa03_sr_6 ) , .B( sa13_sr_6 ) );
  INV_X1 U581 (.ZN( n352 ) , .A( sa03_sr_5 ) );
  XOR2_X1 U582 (.A( n13 ) , .Z( n427 ) , .B( w3_6 ) );
  XOR2_X1 U593 (.Z( N390 ) , .B( sa01_sr_3 ) , .A( w1_27 ) );
  OAI22_X1 U594 (.ZN( N39 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n432 ) , .B1( n433 ) );
  XOR2_X1 U597 (.Z( n436 ) , .B( sa33_sr_4 ) , .A( w3_5 ) );
  XOR2_X1 U598 (.B( n296 ) , .A( n360 ) , .Z( n434 ) );
  XOR2_X1 U599 (.Z( n296 ) , .A( sa03_sr_5 ) , .B( sa13_sr_5 ) );
  INV_X1 U600 (.ZN( n360 ) , .A( sa03_sr_4 ) );
  XOR2_X1 U601 (.A( n11 ) , .Z( n432 ) , .B( w3_5 ) );
  XOR2_X1 U604 (.Z( N388 ) , .B( sa01_sr_5 ) , .A( w1_29 ) );
  OAI22_X1 U613 (.ZN( N38 ) , .A1( n1214 ) , .B2( n1221 ) , .A2( n437 ) , .B1( n438 ) );
  XOR2_X1 U614 (.Z( n438 ) , .A( n439 ) , .B( n440 ) );
  XOR2_X1 U615 (.Z( n440 ) , .B( n441 ) , .A( sa23_sr_4 ) );
  XOR2_X1 U616 (.Z( n441 ) , .B( sa33_sr_3 ) , .A( w3_4 ) );
  XOR2_X1 U617 (.Z( n439 ) , .A( n442 ) , .B( n443 ) );
  XOR2_X1 U618 (.B( n302 ) , .A( n367 ) , .Z( n442 ) );
  XOR2_X1 U619 (.Z( n302 ) , .A( sa03_sr_4 ) , .B( sa13_sr_4 ) );
  INV_X1 U620 (.ZN( n367 ) , .A( sa03_sr_3 ) );
  XOR2_X1 U621 (.Z( n437 ) , .A( n9 ) , .B( w3_4 ) );
  OAI22_X1 U625 (.ZN( N37 ) , .B2( n1114 ) , .A1( n1214 ) , .A2( n444 ) , .B1( n445 ) );
  XOR2_X1 U628 (.Z( n448 ) , .B( sa33_sr_2 ) , .A( w3_3 ) );
  XOR2_X1 U629 (.B( n443 ) , .Z( n446 ) , .A( n449 ) );
  XOR2_X1 U630 (.B( n308 ) , .A( n373 ) , .Z( n449 ) );
  XOR2_X1 U631 (.Z( n308 ) , .A( sa03_sr_3 ) , .B( sa13_sr_3 ) );
  INV_X1 U632 (.ZN( n373 ) , .A( sa03_sr_2 ) );
  XOR2_X1 U633 (.Z( n444 ) , .A( n7 ) , .B( w3_3 ) );
  OAI22_X1 U635 (.ZN( N36 ) , .A1( n1214 ) , .B2( n1220 ) , .A2( n450 ) , .B1( n451 ) );
  XOR2_X1 U636 (.Z( n451 ) , .A( n452 ) , .B( n453 ) );
  XOR2_X1 U637 (.Z( n453 ) , .B( n454 ) , .A( sa23_sr_2 ) );
  XOR2_X1 U638 (.Z( n454 ) , .B( sa33_sr_1 ) , .A( w3_2 ) );
  XOR2_X1 U639 (.B( n316 ) , .A( n380 ) , .Z( n452 ) );
  XOR2_X1 U640 (.Z( n316 ) , .A( sa03_sr_2 ) , .B( sa13_sr_2 ) );
  INV_X1 U641 (.ZN( n380 ) , .A( sa03_sr_1 ) );
  XOR2_X1 U642 (.Z( n450 ) , .A( n5 ) , .B( w3_2 ) );
  OAI22_X1 U644 (.ZN( N35 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n455 ) , .B1( n456 ) );
  XOR2_X1 U647 (.Z( n459 ) , .B( sa33_sr_0 ) , .A( w3_1 ) );
  XOR2_X1 U648 (.B( n443 ) , .Z( n457 ) , .A( n460 ) );
  XOR2_X1 U649 (.B( n323 ) , .A( n386 ) , .Z( n460 ) );
  XOR2_X1 U650 (.Z( n323 ) , .A( sa03_sr_1 ) , .B( sa13_sr_1 ) );
  INV_X1 U651 (.ZN( n386 ) , .A( sa03_sr_0 ) );
  XOR2_X1 U652 (.A( n3 ) , .Z( n455 ) , .B( w3_1 ) );
  OAI22_X1 U654 (.ZN( N34 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n461 ) , .B1( n462 ) );
  XOR2_X1 U656 (.A( n329 ) , .B( n443 ) , .Z( n464 ) );
  XOR2_X1 U657 (.Z( n443 ) , .A( sa03_sr_7 ) , .B( sa33_sr_7 ) );
  XOR2_X1 U658 (.Z( n329 ) , .A( sa03_sr_0 ) , .B( sa13_sr_0 ) );
  XOR2_X1 U660 (.A( n1 ) , .Z( n461 ) , .B( w3_0 ) );
  OAI22_X1 U902 (.ZN( N217 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n639 ) , .B1( n640 ) );
  XOR2_X1 U904 (.Z( n642 ) , .A( n643 ) , .B( n644 ) );
  INV_X1 U906 (.ZN( n645 ) , .A( sa11_sr_7 ) );
  XOR2_X1 U907 (.A( n191 ) , .Z( n639 ) , .B( w1_31 ) );
  OAI22_X1 U909 (.ZN( N216 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n646 ) , .B1( n647 ) );
  XOR2_X1 U911 (.Z( n649 ) , .A( n650 ) , .B( n651 ) );
  XOR2_X1 U913 (.A( n189 ) , .Z( n646 ) , .B( w1_30 ) );
  OAI22_X1 U915 (.ZN( N215 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n652 ) , .B1( n653 ) );
  XOR2_X1 U917 (.Z( n655 ) , .A( n656 ) , .B( n657 ) );
  XOR2_X1 U919 (.A( n187 ) , .Z( n652 ) , .B( w1_29 ) );
  OAI22_X1 U921 (.ZN( N214 ) , .A1( n1109 ) , .B2( n1218 ) , .A2( n658 ) , .B1( n659 ) );
  XOR2_X1 U922 (.Z( n659 ) , .A( n660 ) , .B( n661 ) );
  XOR2_X1 U923 (.Z( n661 ) , .A( n662 ) , .B( n663 ) );
  XOR2_X1 U924 (.Z( n660 ) , .A( n664 ) , .B( n665 ) );
  XNOR2_X1 U925 (.ZN( n664 ) , .B( sa11_sr_4 ) , .A( w1_28 ) );
  XOR2_X1 U926 (.A( n185 ) , .Z( n658 ) , .B( w1_28 ) );
  OAI22_X1 U928 (.ZN( N213 ) , .A1( n1213 ) , .B2( n1218 ) , .A2( n666 ) , .B1( n667 ) );
  XOR2_X1 U930 (.Z( n669 ) , .A( n670 ) , .B( n671 ) );
  XNOR2_X1 U932 (.ZN( n672 ) , .B( sa11_sr_3 ) , .A( w1_27 ) );
  XOR2_X1 U933 (.A( n183 ) , .Z( n666 ) , .B( w1_27 ) );
  OAI22_X1 U935 (.ZN( N212 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n673 ) , .B1( n674 ) );
  XOR2_X1 U937 (.Z( n676 ) , .A( n677 ) , .B( n678 ) );
  XOR2_X1 U939 (.A( n181 ) , .Z( n673 ) , .B( w1_26 ) );
  OAI22_X1 U941 (.ZN( N211 ) , .A1( n1214 ) , .B2( n1218 ) , .A2( n679 ) , .B1( n680 ) );
  XOR2_X1 U943 (.Z( n682 ) , .A( n683 ) , .B( n684 ) );
  XNOR2_X1 U945 (.ZN( n685 ) , .B( sa11_sr_1 ) , .A( w1_25 ) );
  XOR2_X1 U946 (.A( n179 ) , .Z( n679 ) , .B( w1_25 ) );
  OAI22_X1 U948 (.ZN( N210 ) , .A1( n1109 ) , .B2( n1219 ) , .A2( n686 ) , .B1( n687 ) );
  XOR2_X1 U950 (.A( n665 ) , .Z( n689 ) , .B( n690 ) );
  XOR2_X1 U952 (.A( n177 ) , .Z( n686 ) , .B( w1_24 ) );
  OAI22_X1 U954 (.ZN( N201 ) , .A1( n1214 ) , .B2( n1217 ) , .A2( n691 ) , .B1( n692 ) );
  XOR2_X1 U955 (.Z( n692 ) , .A( n693 ) , .B( n694 ) );
  XOR2_X1 U956 (.B( n643 ) , .Z( n694 ) , .A( sa01_sr_7 ) );
  XOR2_X1 U959 (.A( n175 ) , .Z( n691 ) , .B( w1_23 ) );
  OAI22_X1 U961 (.ZN( N200 ) , .A1( n1212 ) , .B2( n1219 ) , .A2( n696 ) , .B1( n697 ) );
  XOR2_X1 U964 (.Z( n700 ) , .B( sa21_sr_5 ) , .A( w1_22 ) );
  XOR2_X1 U967 (.A( n173 ) , .Z( n696 ) , .B( w1_22 ) );
  OAI22_X1 U969 (.ZN( N199 ) , .A1( n1215 ) , .B2( n1218 ) , .A2( n702 ) , .B1( n703 ) );
  XOR2_X1 U970 (.Z( n703 ) , .A( n704 ) , .B( n705 ) );
  XOR2_X1 U971 (.Z( n705 ) , .B( n706 ) , .A( sa11_sr_4 ) );
  XOR2_X1 U972 (.Z( n706 ) , .B( sa21_sr_4 ) , .A( w1_21 ) );
  XNOR2_X1 U973 (.B( n656 ) , .ZN( n704 ) , .A( sa01_sr_5 ) );
  XOR2_X1 U974 (.A( n171 ) , .Z( n702 ) , .B( w1_21 ) );
  OAI22_X1 U976 (.ZN( N198 ) , .A1( n1216 ) , .B2( n1217 ) , .A2( n707 ) , .B1( n708 ) );
  XOR2_X1 U977 (.Z( n708 ) , .A( n709 ) , .B( n710 ) );
  XOR2_X1 U978 (.Z( n710 ) , .B( n711 ) , .A( sa11_sr_3 ) );
  XOR2_X1 U979 (.Z( n711 ) , .B( sa21_sr_3 ) , .A( w1_20 ) );
  XOR2_X1 U980 (.Z( n709 ) , .A( n712 ) , .B( n713 ) );
  XNOR2_X1 U981 (.B( n663 ) , .ZN( n712 ) , .A( sa01_sr_4 ) );
  XOR2_X1 U982 (.A( n169 ) , .Z( n707 ) , .B( w1_20 ) );
  OAI22_X1 U984 (.ZN( N197 ) , .A1( n1109 ) , .B2( n1220 ) , .A2( n714 ) , .B1( n715 ) );
  XOR2_X1 U987 (.Z( n718 ) , .B( sa21_sr_2 ) , .A( w1_19 ) );
  XOR2_X1 U988 (.B( n713 ) , .Z( n716 ) , .A( n719 ) );
  XNOR2_X1 U989 (.B( n670 ) , .ZN( n719 ) , .A( sa01_sr_3 ) );
  XOR2_X1 U990 (.A( n167 ) , .Z( n714 ) , .B( w1_19 ) );
  OAI22_X1 U992 (.ZN( N196 ) , .A1( n1212 ) , .B2( n1218 ) , .A2( n720 ) , .B1( n721 ) );
  XOR2_X1 U995 (.Z( n724 ) , .B( sa21_sr_1 ) , .A( w1_18 ) );
  XNOR2_X1 U996 (.B( n677 ) , .ZN( n722 ) , .A( sa01_sr_2 ) );
  XOR2_X1 U997 (.A( n165 ) , .Z( n720 ) , .B( w1_18 ) );
  OAI22_X1 U999 (.ZN( N195 ) , .A1( n1215 ) , .B2( n1221 ) , .A2( n725 ) , .B1( n726 ) );
  INV_X1 u0_U203 (.A( u0_n250 ) , .ZN( w3_13 ) );
  INV_X1 u0_U206 (.A( u0_n254 ) , .ZN( w3_14 ) );
  INV_X1 u0_U210 (.A( u0_n258 ) , .ZN( w3_12 ) );
  INV_X1 u0_U230 (.A( u0_n264 ) , .ZN( w3_15 ) );
  XOR2_X1 u0_U294 (.Z( u0_n74 ) , .A( u0_n76 ) , .B( w3_28 ) );
  XOR2_X1 u0_U297 (.Z( u0_n83 ) , .A( u0_n85 ) , .B( w3_25 ) );
  XOR2_X1 u0_U307 (.Z( u0_n113 ) , .A( u0_n115 ) , .B( w3_15 ) );
  XOR2_X1 u0_U308 (.Z( u0_n116 ) , .A( u0_n118 ) , .B( w3_14 ) );
  XOR2_X1 u0_U309 (.Z( u0_n119 ) , .A( u0_n121 ) , .B( w3_13 ) );
  XOR2_X1 u0_U310 (.Z( u0_n122 ) , .A( u0_n124 ) , .B( w3_12 ) );
  XOR2_X1 u0_U312 (.Z( u0_n128 ) , .A( u0_n130 ) , .B( w3_10 ) );
  XOR2_X1 u0_U326 (.A( u0_n168 ) , .Z( u0_n76 ) , .B( w2_28 ) );
  XOR2_X1 u0_U329 (.A( u0_n174 ) , .Z( u0_n85 ) , .B( w2_25 ) );
  XOR2_X1 u0_U339 (.Z( u0_n115 ) , .A( u0_n194 ) , .B( w2_15 ) );
  XOR2_X1 u0_U340 (.Z( u0_n118 ) , .A( u0_n196 ) , .B( w2_14 ) );
  XOR2_X1 u0_U341 (.Z( u0_n121 ) , .A( u0_n198 ) , .B( w2_13 ) );
  XOR2_X1 u0_U342 (.Z( u0_n124 ) , .A( u0_n200 ) , .B( w2_12 ) );
  XOR2_X1 u0_U344 (.Z( u0_n130 ) , .A( u0_n204 ) , .B( w2_10 ) );
  XOR2_X1 u0_U361 (.Z( u0_n168 ) , .A( u0_n7 ) , .B( w1_28 ) );
  XOR2_X1 u0_U367 (.A( u0_n13 ) , .Z( u0_n174 ) , .B( w1_25 ) );
  XOR2_X1 u0_U387 (.Z( u0_n194 ) , .A( u0_n33 ) , .B( w1_15 ) );
  XOR2_X1 u0_U389 (.Z( u0_n196 ) , .A( u0_n35 ) , .B( w1_14 ) );
  XOR2_X1 u0_U391 (.Z( u0_n198 ) , .A( u0_n37 ) , .B( w1_13 ) );
  XOR2_X1 u0_U393 (.Z( u0_n200 ) , .A( u0_n39 ) , .B( w1_12 ) );
  XOR2_X1 u0_U397 (.Z( u0_n204 ) , .A( u0_n43 ) , .B( w1_10 ) );
endmodule

