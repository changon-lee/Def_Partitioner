module aes_aes ( clk, key, ld, rst, text_in, done, text_out );
  input clk;
  input [127:0] key;
  input ld;
  input rst;
  input [127:0] text_in;
  output done;
  output [127:0] text_out;

  wire sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, 
       sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, sa01_0, 
       sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa01_sr_0, sa01_sr_1, 
       sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_0, sa02_1, sa02_2, 
       sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, 
       sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa03_0, sa03_1, sa03_2, sa03_3, sa03_4, 
       sa03_5, sa03_6, sa03_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, 
       sa03_sr_6, sa03_sr_7, sa10_0, sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, 
       sa10_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, 
       sa11_0, sa11_1, sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa11_sr_0, 
       sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa12_0, sa12_1, 
       sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, 
       sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, sa13_0, sa13_1, sa13_2, sa13_3, 
       sa13_4, sa13_5, sa13_6, sa13_7, sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, 
       sa13_sr_5, sa13_sr_6, sa13_sr_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, 
       sa20_6, sa20_7, sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, 
       sa21_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, sa21_sr_7, 
       sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa23_0, 
       sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa23_sr_0, sa23_sr_1, 
       sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa30_0, sa30_1, sa30_2, 
       sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa30_sr_0, sa30_sr_1, sa30_sr_2, sa30_sr_3, 
       sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, sa31_0, sa31_1, sa31_2, sa31_3, sa31_4, 
       sa31_5, sa31_6, sa31_7, sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, 
       sa31_sr_6, sa31_sr_7, sa32_0, sa32_1, sa32_2, sa32_3, sa32_4, sa32_5, sa32_6, 
       sa32_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, 
       sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, sa33_5, sa33_6, sa33_7, sa33_sr_0, 
       sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_n268, u0_n270, 
       u0_n272, u0_n274, u0_subword_0, u0_subword_1, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, u0_subword_14, 
       u0_subword_15, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_2, u0_subword_20, u0_subword_21, u0_subword_22, 
       u0_subword_23, u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7, u0_subword_8, u0_subword_9, w3_0, 
       w3_1, w3_10, w3_11, w3_2, w3_24, w3_25, w3_26, w3_27, w3_28, 
       w3_29, w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, 
       w3_9 ;

  aes_aes_die_0 u0 ( clk, key, ld, rst, text_in, done, text_out, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, sa00_sr_6, sa00_sr_7, 
      sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, 
      sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa03_sr_0, sa03_sr_1, 
      sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, 
      sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, sa10_sr_7, sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, 
      sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, 
      sa12_sr_5, sa12_sr_6, sa12_sr_7, sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, 
      sa13_sr_6, sa13_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, 
      sa21_sr_7, sa22_sr_0, sa22_sr_1, sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, 
      sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, sa30_sr_0, 
      sa30_sr_1, sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7, sa31_sr_0, sa31_sr_1, 
      sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, 
      sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, sa33_sr_0, sa33_sr_1, sa33_sr_2, sa33_sr_3, 
      sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_subword_0, u0_subword_1, u0_subword_10, u0_subword_11, u0_subword_12, 
      u0_subword_13, u0_subword_14, u0_subword_15, u0_subword_16, u0_subword_17, u0_subword_18, u0_subword_19, u0_subword_2, u0_subword_20, 
      u0_subword_21, u0_subword_22, u0_subword_23, u0_subword_3, u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7, u0_subword_8, 
      u0_subword_9, sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, 
      sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, 
      sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa03_0, sa03_1, 
      sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa10_0, sa10_1, sa10_2, 
      sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, sa11_2, sa11_3, 
      sa11_4, sa11_5, sa11_6, sa11_7, sa12_0, sa12_1, sa12_2, sa12_3, sa12_4, 
      sa12_5, sa12_6, sa12_7, sa13_0, sa13_1, sa13_2, sa13_3, sa13_4, sa13_5, 
      sa13_6, sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, sa20_4, sa20_5, sa20_6, 
      sa20_7, sa21_0, sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, 
      sa23_0, sa23_1, sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, 
      sa30_1, sa30_2, sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa31_0, sa31_1, 
      sa31_2, sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, sa32_0, sa32_1, sa32_2, 
      sa32_3, sa32_4, sa32_5, sa32_6, sa32_7, sa33_0, sa33_1, sa33_2, sa33_3, 
      sa33_4, sa33_5, sa33_6, sa33_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_0, 
      w3_1, w3_10, w3_11, w3_2, w3_24, w3_25, w3_26, w3_27, w3_28, 
      w3_29, w3_3, w3_30, w3_31, w3_4, w3_5, w3_6, w3_7, w3_8, 
      w3_9 );
  aes_aes_die_1 u1 ( sa00_0, sa00_1, sa00_2, sa00_3, sa00_4, sa00_5, sa00_6, sa00_7, sa03_0, 
      sa03_1, sa03_2, sa03_3, sa03_4, sa03_5, sa03_6, sa03_7, sa12_0, sa12_1, 
      sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa31_0, sa31_1, sa31_2, 
      sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, w3_0, w3_1, w3_2, w3_24, 
      w3_25, w3_26, w3_27, w3_28, w3_29, w3_3, w3_30, w3_31, w3_4, 
      w3_5, w3_6, w3_7, sa00_sr_0, sa00_sr_1, sa00_sr_2, sa00_sr_3, sa00_sr_4, sa00_sr_5, 
      sa00_sr_6, sa00_sr_7, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, 
      sa03_sr_7, sa11_sr_0, sa11_sr_1, sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, 
      sa32_sr_0, sa32_sr_1, sa32_sr_2, sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, u0_subword_0, 
      u0_subword_1, u0_subword_10, u0_subword_11, u0_subword_12, u0_subword_13, u0_subword_14, u0_subword_15, u0_subword_2, u0_subword_3, 
      u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7, u0_subword_8, u0_subword_9 );
  aes_aes_die_2 u2 ( sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa10_0, 
      sa10_1, sa10_2, sa10_3, sa10_4, sa10_5, sa10_6, sa10_7, sa11_0, sa11_1, 
      sa11_2, sa11_3, sa11_4, sa11_5, sa11_6, sa11_7, sa13_0, sa13_1, sa13_2, 
      sa13_3, sa13_4, sa13_5, sa13_6, sa13_7, sa20_0, sa20_1, sa20_2, sa20_3, 
      sa20_4, sa20_5, sa20_6, sa20_7, sa33_0, sa33_1, sa33_2, sa33_3, sa33_4, 
      sa33_5, sa33_6, sa33_7, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, 
      sa01_sr_6, sa01_sr_7, sa10_sr_0, sa10_sr_1, sa10_sr_2, sa10_sr_3, sa10_sr_4, sa10_sr_5, sa10_sr_6, 
      sa10_sr_7, sa12_sr_0, sa12_sr_1, sa12_sr_2, sa12_sr_3, sa12_sr_4, sa12_sr_5, sa12_sr_6, sa12_sr_7, 
      sa13_sr_0, sa13_sr_1, sa13_sr_2, sa13_sr_3, sa13_sr_4, sa13_sr_5, sa13_sr_6, sa13_sr_7, sa22_sr_0, 
      sa22_sr_1, sa22_sr_2, sa22_sr_3, sa22_sr_4, sa22_sr_5, sa22_sr_6, sa22_sr_7, sa30_sr_0, sa30_sr_1, 
      sa30_sr_2, sa30_sr_3, sa30_sr_4, sa30_sr_5, sa30_sr_6, sa30_sr_7 );
  aes_aes_die_3 u3 ( sa02_0, sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa21_0, 
      sa21_1, sa21_2, sa21_3, sa21_4, sa21_5, sa21_6, sa21_7, sa23_0, sa23_1, 
      sa23_2, sa23_3, sa23_4, sa23_5, sa23_6, sa23_7, sa30_0, sa30_1, sa30_2, 
      sa30_3, sa30_4, sa30_5, sa30_6, sa30_7, sa32_0, sa32_1, sa32_2, sa32_3, 
      sa32_4, sa32_5, sa32_6, sa32_7, u0_n268, u0_n270, u0_n272, u0_n274, w3_10, 
      w3_11, w3_8, w3_9, sa02_sr_0, sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, 
      sa02_sr_6, sa02_sr_7, sa21_sr_0, sa21_sr_1, sa21_sr_2, sa21_sr_3, sa21_sr_4, sa21_sr_5, sa21_sr_6, 
      sa21_sr_7, sa23_sr_0, sa23_sr_1, sa23_sr_2, sa23_sr_3, sa23_sr_4, sa23_sr_5, sa23_sr_6, sa23_sr_7, 
      sa31_sr_0, sa31_sr_1, sa31_sr_2, sa31_sr_3, sa31_sr_4, sa31_sr_5, sa31_sr_6, sa31_sr_7, sa33_sr_0, 
      sa33_sr_1, sa33_sr_2, sa33_sr_3, sa33_sr_4, sa33_sr_5, sa33_sr_6, sa33_sr_7, u0_subword_16, u0_subword_17, 
      u0_subword_18, u0_subword_19, u0_subword_20, u0_subword_21, u0_subword_22, u0_subword_23 );
endmodule
