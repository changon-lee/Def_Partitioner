module des_des_die_5 ( u1_L0_12, u1_L0_14, u1_L0_22, u1_L0_25, u1_L0_3, u1_L0_32, u1_L0_7, u1_L0_8, u1_L11_12, 
       u1_L11_15, u1_L11_16, u1_L11_21, u1_L11_22, u1_L11_24, u1_L11_27, u1_L11_30, u1_L11_32, u1_L11_5, 
       u1_L11_6, u1_L11_7, u1_L12_11, u1_L12_14, u1_L12_19, u1_L12_25, u1_L12_29, u1_L12_3, u1_L12_4, 
       u1_L12_8, u1_L1_1, u1_L1_10, u1_L1_13, u1_L1_16, u1_L1_17, u1_L1_18, u1_L1_2, u1_L1_20, 
       u1_L1_23, u1_L1_24, u1_L1_26, u1_L1_28, u1_L1_30, u1_L1_31, u1_L1_6, u1_L1_9, u1_L3_16, 
       u1_L3_17, u1_L3_23, u1_L3_24, u1_L3_30, u1_L3_31, u1_L3_6, u1_L3_9, u1_L5_11, u1_L5_17, 
       u1_L5_19, u1_L5_23, u1_L5_29, u1_L5_31, u1_L5_4, u1_L5_9, u1_L6_11, u1_L6_14, u1_L6_19, 
       u1_L6_25, u1_L6_29, u1_L6_3, u1_L6_4, u1_L6_8, u1_L7_14, u1_L7_25, u1_L7_3, u1_L7_8, 
       u1_L8_14, u1_L8_25, u1_L8_3, u1_L8_8, u1_R0_16, u1_R0_17, u1_R0_18, u1_R0_19, u1_R0_20, 
       u1_R0_21, u1_R0_24, u1_R0_25, u1_R0_26, u1_R0_27, u1_R0_28, u1_R0_29, u1_R11_1, u1_R11_10, 
       u1_R11_11, u1_R11_12, u1_R11_13, u1_R11_24, u1_R11_25, u1_R11_26, u1_R11_27, u1_R11_28, u1_R11_29, 
       u1_R11_30, u1_R11_31, u1_R11_32, u1_R11_8, u1_R11_9, u1_R12_16, u1_R12_17, u1_R12_18, u1_R12_19, 
       u1_R12_20, u1_R12_21, u1_R12_22, u1_R12_23, u1_R12_24, u1_R12_25, u1_R1_1, u1_R1_10, u1_R1_11, 
       u1_R1_12, u1_R1_13, u1_R1_14, u1_R1_15, u1_R1_16, u1_R1_17, u1_R1_2, u1_R1_3, u1_R1_32, 
       u1_R1_4, u1_R1_5, u1_R1_6, u1_R1_7, u1_R1_8, u1_R1_9, u1_R3_1, u1_R3_10, u1_R3_11, 
       u1_R3_12, u1_R3_13, u1_R3_2, u1_R3_3, u1_R3_32, u1_R3_4, u1_R3_5, u1_R3_8, u1_R3_9, 
       u1_R5_1, u1_R5_2, u1_R5_20, u1_R5_21, u1_R5_22, u1_R5_23, u1_R5_24, u1_R5_25, u1_R5_3, 
       u1_R5_32, u1_R5_4, u1_R5_5, u1_R6_16, u1_R6_17, u1_R6_18, u1_R6_19, u1_R6_20, u1_R6_21, 
       u1_R6_22, u1_R6_23, u1_R6_24, u1_R6_25, u1_R7_16, u1_R7_17, u1_R7_18, u1_R7_19, u1_R7_20, 
       u1_R7_21, u1_R8_16, u1_R8_17, u1_R8_18, u1_R8_19, u1_R8_20, u1_R8_21, u1_uk_K_r0_15, u1_uk_K_r0_22, 
       u1_uk_K_r0_28, u1_uk_K_r0_49, u1_uk_K_r0_7, u1_uk_K_r11_11, u1_uk_K_r11_20, u1_uk_K_r11_27, u1_uk_K_r11_29, u1_uk_K_r11_48, u1_uk_K_r11_6, 
       u1_uk_K_r11_8, u1_uk_K_r12_1, u1_uk_K_r12_30, u1_uk_K_r12_36, u1_uk_K_r12_42, u1_uk_K_r12_44, u1_uk_K_r12_7, u1_uk_K_r1_10, u1_uk_K_r1_17, 
       u1_uk_K_r1_18, u1_uk_K_r1_33, u1_uk_K_r1_41, u1_uk_K_r1_47, u1_uk_K_r1_6, u1_uk_K_r3_10, u1_uk_K_r3_34, u1_uk_K_r3_4, u1_uk_K_r5_0, 
       u1_uk_K_r5_1, u1_uk_K_r5_10, u1_uk_K_r5_16, u1_uk_K_r5_21, u1_uk_K_r5_35, u1_uk_K_r5_37, u1_uk_K_r5_39, u1_uk_K_r5_4, u1_uk_K_r5_41, 
       u1_uk_K_r5_51, u1_uk_K_r6_14, u1_uk_K_r6_21, u1_uk_K_r6_28, u1_uk_K_r6_29, u1_uk_K_r6_35, u1_uk_K_r6_51, u1_uk_K_r7_15, u1_uk_K_r7_2, 
       u1_uk_K_r7_29, u1_uk_K_r7_8, u1_uk_K_r7_9, u1_uk_K_r8_43, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n110, u1_uk_n117, 
       u1_uk_n118, u1_uk_n1260, u1_uk_n1265, u1_uk_n1266, u1_uk_n1267, u1_uk_n1276, u1_uk_n128, u1_uk_n1281, u1_uk_n1282, 
       u1_uk_n1289, u1_uk_n129, u1_uk_n1294, u1_uk_n1295, u1_uk_n1296, u1_uk_n1304, u1_uk_n1310, u1_uk_n1311, u1_uk_n1312, 
       u1_uk_n1315, u1_uk_n1316, u1_uk_n1317, u1_uk_n1319, u1_uk_n1320, u1_uk_n1321, u1_uk_n1323, u1_uk_n1324, u1_uk_n1325, 
       u1_uk_n1326, u1_uk_n1331, u1_uk_n1332, u1_uk_n1336, u1_uk_n1340, u1_uk_n1341, u1_uk_n1346, u1_uk_n1347, u1_uk_n1348, 
       u1_uk_n1397, u1_uk_n1398, u1_uk_n1399, u1_uk_n1402, u1_uk_n1403, u1_uk_n1404, u1_uk_n1405, u1_uk_n1409, u1_uk_n1410, 
       u1_uk_n1411, u1_uk_n1417, u1_uk_n142, u1_uk_n1422, u1_uk_n1424, u1_uk_n1429, u1_uk_n1436, u1_uk_n146, u1_uk_n1482, 
       u1_uk_n1484, u1_uk_n1487, u1_uk_n1492, u1_uk_n1494, u1_uk_n1495, u1_uk_n1504, u1_uk_n1508, u1_uk_n1514, u1_uk_n1517, 
       u1_uk_n1527, u1_uk_n1528, u1_uk_n1529, u1_uk_n1533, u1_uk_n1534, u1_uk_n1540, u1_uk_n1541, u1_uk_n1547, u1_uk_n1554, 
       u1_uk_n1555, u1_uk_n1556, u1_uk_n1560, u1_uk_n1562, u1_uk_n1563, u1_uk_n1567, u1_uk_n1568, u1_uk_n1595, u1_uk_n1599, 
       u1_uk_n1600, u1_uk_n1607, u1_uk_n1608, u1_uk_n161, u1_uk_n1614, u1_uk_n1615, u1_uk_n1623, u1_uk_n1627, u1_uk_n1628, 
       u1_uk_n1632, u1_uk_n1639, u1_uk_n164, u1_uk_n1640, u1_uk_n1641, u1_uk_n1647, u1_uk_n1655, u1_uk_n1656, u1_uk_n1753, 
       u1_uk_n1754, u1_uk_n1755, u1_uk_n1756, u1_uk_n1761, u1_uk_n1763, u1_uk_n1764, u1_uk_n1766, u1_uk_n1768, u1_uk_n1769, 
       u1_uk_n1773, u1_uk_n1774, u1_uk_n1775, u1_uk_n1776, u1_uk_n1780, u1_uk_n1782, u1_uk_n1784, u1_uk_n1785, u1_uk_n1791, 
       u1_uk_n1792, u1_uk_n1793, u1_uk_n1799, u1_uk_n1800, u1_uk_n1806, u1_uk_n1811, u1_uk_n1815, u1_uk_n182, u1_uk_n1821, 
       u1_uk_n1822, u1_uk_n1827, u1_uk_n1833, u1_uk_n1837, u1_uk_n1838, u1_uk_n1839, u1_uk_n187, u1_uk_n188, u1_uk_n203, 
       u1_uk_n207, u1_uk_n230, u1_uk_n231, u1_uk_n250, u1_uk_n251, u1_uk_n252, u1_uk_n257, u1_uk_n291, u1_uk_n294, 
       u1_uk_n297, u1_uk_n298, u1_uk_n60, u1_uk_n63, u1_uk_n83, u1_uk_n92, u1_uk_n94, u2_FP_33, u2_FP_60, 
       u2_FP_61, u2_FP_62, u2_FP_63, u2_FP_64, u2_K16_44, u2_K16_47, u2_L14_15, u2_L14_21, u2_L14_27, 
       u2_L14_5, u2_L5_1, u2_L5_10, u2_L5_20, u2_L5_26, u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_15, 
       u2_R5_16, u2_R5_17, u2_uk_K_r14_16, u2_uk_K_r14_9, u2_uk_K_r5_18, u2_uk_K_r5_19, u2_uk_K_r5_40, u2_uk_n100, u2_uk_n1079, 
       u2_uk_n1081, u2_uk_n1082, u2_uk_n11, u2_uk_n118, u2_uk_n1189, u2_uk_n1200, u2_uk_n1208, u2_uk_n1217, u2_uk_n1220, 
       u2_uk_n1223, u2_uk_n128, u2_uk_n129, u2_uk_n1453, u2_uk_n1465, u2_uk_n1468, u2_uk_n1475, u2_uk_n1496, u2_uk_n161, 
       u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n217, u2_uk_n231, u2_uk_n238, u2_uk_n31, u2_uk_n94, u1_N133, u1_N136, u1_N143, u1_N144, u1_N150, u1_N151, u1_N157, u1_N158, u1_N195, 
        u1_N200, u1_N202, u1_N208, u1_N210, u1_N214, u1_N220, u1_N222, u1_N226, u1_N227, 
        u1_N231, u1_N234, u1_N237, u1_N242, u1_N248, u1_N252, u1_N258, u1_N263, u1_N269, 
        u1_N280, u1_N290, u1_N295, u1_N301, u1_N312, u1_N34, u1_N38, u1_N388, u1_N389, 
        u1_N39, u1_N390, u1_N395, u1_N398, u1_N399, u1_N404, u1_N405, u1_N407, u1_N410, 
        u1_N413, u1_N415, u1_N418, u1_N419, u1_N423, u1_N426, u1_N429, u1_N43, u1_N434, 
        u1_N440, u1_N444, u1_N45, u1_N53, u1_N56, u1_N63, u1_N64, u1_N65, u1_N69, 
        u1_N72, u1_N73, u1_N76, u1_N79, u1_N80, u1_N81, u1_N83, u1_N86, u1_N87, 
        u1_N89, u1_N91, u1_N93, u1_N94, u1_uk_n10, u1_uk_n11, u1_uk_n141, u1_uk_n145, u1_uk_n147, 
        u1_uk_n148, u1_uk_n155, u1_uk_n162, u1_uk_n163, u1_uk_n17, u1_uk_n191, u1_uk_n202, u1_uk_n208, u1_uk_n209, 
        u1_uk_n214, u1_uk_n217, u1_uk_n220, u1_uk_n222, u1_uk_n223, u1_uk_n238, u1_uk_n240, u1_uk_n242, u1_uk_n27, 
        u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n286, u1_uk_n292, u1_uk_n31, u1_uk_n93, u1_uk_n99, u2_FP_15, 
        u2_FP_21, u2_FP_27, u2_FP_5, u2_N192, u2_N201, u2_N211, u2_N217 );
  input u1_L0_12, u1_L0_14, u1_L0_22, u1_L0_25, u1_L0_3, u1_L0_32, u1_L0_7, u1_L0_8, u1_L11_12, 
        u1_L11_15, u1_L11_16, u1_L11_21, u1_L11_22, u1_L11_24, u1_L11_27, u1_L11_30, u1_L11_32, u1_L11_5, 
        u1_L11_6, u1_L11_7, u1_L12_11, u1_L12_14, u1_L12_19, u1_L12_25, u1_L12_29, u1_L12_3, u1_L12_4, 
        u1_L12_8, u1_L1_1, u1_L1_10, u1_L1_13, u1_L1_16, u1_L1_17, u1_L1_18, u1_L1_2, u1_L1_20, 
        u1_L1_23, u1_L1_24, u1_L1_26, u1_L1_28, u1_L1_30, u1_L1_31, u1_L1_6, u1_L1_9, u1_L3_16, 
        u1_L3_17, u1_L3_23, u1_L3_24, u1_L3_30, u1_L3_31, u1_L3_6, u1_L3_9, u1_L5_11, u1_L5_17, 
        u1_L5_19, u1_L5_23, u1_L5_29, u1_L5_31, u1_L5_4, u1_L5_9, u1_L6_11, u1_L6_14, u1_L6_19, 
        u1_L6_25, u1_L6_29, u1_L6_3, u1_L6_4, u1_L6_8, u1_L7_14, u1_L7_25, u1_L7_3, u1_L7_8, 
        u1_L8_14, u1_L8_25, u1_L8_3, u1_L8_8, u1_R0_16, u1_R0_17, u1_R0_18, u1_R0_19, u1_R0_20, 
        u1_R0_21, u1_R0_24, u1_R0_25, u1_R0_26, u1_R0_27, u1_R0_28, u1_R0_29, u1_R11_1, u1_R11_10, 
        u1_R11_11, u1_R11_12, u1_R11_13, u1_R11_24, u1_R11_25, u1_R11_26, u1_R11_27, u1_R11_28, u1_R11_29, 
        u1_R11_30, u1_R11_31, u1_R11_32, u1_R11_8, u1_R11_9, u1_R12_16, u1_R12_17, u1_R12_18, u1_R12_19, 
        u1_R12_20, u1_R12_21, u1_R12_22, u1_R12_23, u1_R12_24, u1_R12_25, u1_R1_1, u1_R1_10, u1_R1_11, 
        u1_R1_12, u1_R1_13, u1_R1_14, u1_R1_15, u1_R1_16, u1_R1_17, u1_R1_2, u1_R1_3, u1_R1_32, 
        u1_R1_4, u1_R1_5, u1_R1_6, u1_R1_7, u1_R1_8, u1_R1_9, u1_R3_1, u1_R3_10, u1_R3_11, 
        u1_R3_12, u1_R3_13, u1_R3_2, u1_R3_3, u1_R3_32, u1_R3_4, u1_R3_5, u1_R3_8, u1_R3_9, 
        u1_R5_1, u1_R5_2, u1_R5_20, u1_R5_21, u1_R5_22, u1_R5_23, u1_R5_24, u1_R5_25, u1_R5_3, 
        u1_R5_32, u1_R5_4, u1_R5_5, u1_R6_16, u1_R6_17, u1_R6_18, u1_R6_19, u1_R6_20, u1_R6_21, 
        u1_R6_22, u1_R6_23, u1_R6_24, u1_R6_25, u1_R7_16, u1_R7_17, u1_R7_18, u1_R7_19, u1_R7_20, 
        u1_R7_21, u1_R8_16, u1_R8_17, u1_R8_18, u1_R8_19, u1_R8_20, u1_R8_21, u1_uk_K_r0_15, u1_uk_K_r0_22, 
        u1_uk_K_r0_28, u1_uk_K_r0_49, u1_uk_K_r0_7, u1_uk_K_r11_11, u1_uk_K_r11_20, u1_uk_K_r11_27, u1_uk_K_r11_29, u1_uk_K_r11_48, u1_uk_K_r11_6, 
        u1_uk_K_r11_8, u1_uk_K_r12_1, u1_uk_K_r12_30, u1_uk_K_r12_36, u1_uk_K_r12_42, u1_uk_K_r12_44, u1_uk_K_r12_7, u1_uk_K_r1_10, u1_uk_K_r1_17, 
        u1_uk_K_r1_18, u1_uk_K_r1_33, u1_uk_K_r1_41, u1_uk_K_r1_47, u1_uk_K_r1_6, u1_uk_K_r3_10, u1_uk_K_r3_34, u1_uk_K_r3_4, u1_uk_K_r5_0, 
        u1_uk_K_r5_1, u1_uk_K_r5_10, u1_uk_K_r5_16, u1_uk_K_r5_21, u1_uk_K_r5_35, u1_uk_K_r5_37, u1_uk_K_r5_39, u1_uk_K_r5_4, u1_uk_K_r5_41, 
        u1_uk_K_r5_51, u1_uk_K_r6_14, u1_uk_K_r6_21, u1_uk_K_r6_28, u1_uk_K_r6_29, u1_uk_K_r6_35, u1_uk_K_r6_51, u1_uk_K_r7_15, u1_uk_K_r7_2, 
        u1_uk_K_r7_29, u1_uk_K_r7_8, u1_uk_K_r7_9, u1_uk_K_r8_43, u1_uk_n100, u1_uk_n102, u1_uk_n109, u1_uk_n110, u1_uk_n117, 
        u1_uk_n118, u1_uk_n1260, u1_uk_n1265, u1_uk_n1266, u1_uk_n1267, u1_uk_n1276, u1_uk_n128, u1_uk_n1281, u1_uk_n1282, 
        u1_uk_n1289, u1_uk_n129, u1_uk_n1294, u1_uk_n1295, u1_uk_n1296, u1_uk_n1304, u1_uk_n1310, u1_uk_n1311, u1_uk_n1312, 
        u1_uk_n1315, u1_uk_n1316, u1_uk_n1317, u1_uk_n1319, u1_uk_n1320, u1_uk_n1321, u1_uk_n1323, u1_uk_n1324, u1_uk_n1325, 
        u1_uk_n1326, u1_uk_n1331, u1_uk_n1332, u1_uk_n1336, u1_uk_n1340, u1_uk_n1341, u1_uk_n1346, u1_uk_n1347, u1_uk_n1348, 
        u1_uk_n1397, u1_uk_n1398, u1_uk_n1399, u1_uk_n1402, u1_uk_n1403, u1_uk_n1404, u1_uk_n1405, u1_uk_n1409, u1_uk_n1410, 
        u1_uk_n1411, u1_uk_n1417, u1_uk_n142, u1_uk_n1422, u1_uk_n1424, u1_uk_n1429, u1_uk_n1436, u1_uk_n146, u1_uk_n1482, 
        u1_uk_n1484, u1_uk_n1487, u1_uk_n1492, u1_uk_n1494, u1_uk_n1495, u1_uk_n1504, u1_uk_n1508, u1_uk_n1514, u1_uk_n1517, 
        u1_uk_n1527, u1_uk_n1528, u1_uk_n1529, u1_uk_n1533, u1_uk_n1534, u1_uk_n1540, u1_uk_n1541, u1_uk_n1547, u1_uk_n1554, 
        u1_uk_n1555, u1_uk_n1556, u1_uk_n1560, u1_uk_n1562, u1_uk_n1563, u1_uk_n1567, u1_uk_n1568, u1_uk_n1595, u1_uk_n1599, 
        u1_uk_n1600, u1_uk_n1607, u1_uk_n1608, u1_uk_n161, u1_uk_n1614, u1_uk_n1615, u1_uk_n1623, u1_uk_n1627, u1_uk_n1628, 
        u1_uk_n1632, u1_uk_n1639, u1_uk_n164, u1_uk_n1640, u1_uk_n1641, u1_uk_n1647, u1_uk_n1655, u1_uk_n1656, u1_uk_n1753, 
        u1_uk_n1754, u1_uk_n1755, u1_uk_n1756, u1_uk_n1761, u1_uk_n1763, u1_uk_n1764, u1_uk_n1766, u1_uk_n1768, u1_uk_n1769, 
        u1_uk_n1773, u1_uk_n1774, u1_uk_n1775, u1_uk_n1776, u1_uk_n1780, u1_uk_n1782, u1_uk_n1784, u1_uk_n1785, u1_uk_n1791, 
        u1_uk_n1792, u1_uk_n1793, u1_uk_n1799, u1_uk_n1800, u1_uk_n1806, u1_uk_n1811, u1_uk_n1815, u1_uk_n182, u1_uk_n1821, 
        u1_uk_n1822, u1_uk_n1827, u1_uk_n1833, u1_uk_n1837, u1_uk_n1838, u1_uk_n1839, u1_uk_n187, u1_uk_n188, u1_uk_n203, 
        u1_uk_n207, u1_uk_n230, u1_uk_n231, u1_uk_n250, u1_uk_n251, u1_uk_n252, u1_uk_n257, u1_uk_n291, u1_uk_n294, 
        u1_uk_n297, u1_uk_n298, u1_uk_n60, u1_uk_n63, u1_uk_n83, u1_uk_n92, u1_uk_n94, u2_FP_33, u2_FP_60, 
        u2_FP_61, u2_FP_62, u2_FP_63, u2_FP_64, u2_K16_44, u2_K16_47, u2_L14_15, u2_L14_21, u2_L14_27, 
        u2_L14_5, u2_L5_1, u2_L5_10, u2_L5_20, u2_L5_26, u2_R5_12, u2_R5_13, u2_R5_14, u2_R5_15, 
        u2_R5_16, u2_R5_17, u2_uk_K_r14_16, u2_uk_K_r14_9, u2_uk_K_r5_18, u2_uk_K_r5_19, u2_uk_K_r5_40, u2_uk_n100, u2_uk_n1079, 
        u2_uk_n1081, u2_uk_n1082, u2_uk_n11, u2_uk_n118, u2_uk_n1189, u2_uk_n1200, u2_uk_n1208, u2_uk_n1217, u2_uk_n1220, 
        u2_uk_n1223, u2_uk_n128, u2_uk_n129, u2_uk_n1453, u2_uk_n1465, u2_uk_n1468, u2_uk_n1475, u2_uk_n1496, u2_uk_n161, 
        u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n217, u2_uk_n231, u2_uk_n238, u2_uk_n31, u2_uk_n94;
  output u1_N133, u1_N136, u1_N143, u1_N144, u1_N150, u1_N151, u1_N157, u1_N158, u1_N195, 
        u1_N200, u1_N202, u1_N208, u1_N210, u1_N214, u1_N220, u1_N222, u1_N226, u1_N227, 
        u1_N231, u1_N234, u1_N237, u1_N242, u1_N248, u1_N252, u1_N258, u1_N263, u1_N269, 
        u1_N280, u1_N290, u1_N295, u1_N301, u1_N312, u1_N34, u1_N38, u1_N388, u1_N389, 
        u1_N39, u1_N390, u1_N395, u1_N398, u1_N399, u1_N404, u1_N405, u1_N407, u1_N410, 
        u1_N413, u1_N415, u1_N418, u1_N419, u1_N423, u1_N426, u1_N429, u1_N43, u1_N434, 
        u1_N440, u1_N444, u1_N45, u1_N53, u1_N56, u1_N63, u1_N64, u1_N65, u1_N69, 
        u1_N72, u1_N73, u1_N76, u1_N79, u1_N80, u1_N81, u1_N83, u1_N86, u1_N87, 
        u1_N89, u1_N91, u1_N93, u1_N94, u1_uk_n10, u1_uk_n11, u1_uk_n141, u1_uk_n145, u1_uk_n147, 
        u1_uk_n148, u1_uk_n155, u1_uk_n162, u1_uk_n163, u1_uk_n17, u1_uk_n191, u1_uk_n202, u1_uk_n208, u1_uk_n209, 
        u1_uk_n214, u1_uk_n217, u1_uk_n220, u1_uk_n222, u1_uk_n223, u1_uk_n238, u1_uk_n240, u1_uk_n242, u1_uk_n27, 
        u1_uk_n271, u1_uk_n277, u1_uk_n279, u1_uk_n286, u1_uk_n292, u1_uk_n31, u1_uk_n93, u1_uk_n99, u2_FP_15, 
        u2_FP_21, u2_FP_27, u2_FP_5, u2_N192, u2_N201, u2_N211, u2_N217;
  wire u1_K10_25, u1_K10_26, u1_K10_27, u1_K10_28, u1_K10_29, u1_K10_30, u1_K13_13, u1_K13_14, u1_K13_15, 
       u1_K13_16, u1_K13_17, u1_K13_18, u1_K13_37, u1_K13_38, u1_K13_39, u1_K13_40, u1_K13_41, u1_K13_42, 
       u1_K13_43, u1_K13_44, u1_K13_45, u1_K13_46, u1_K13_47, u1_K13_48, u1_K14_25, u1_K14_26, u1_K14_27, 
       u1_K14_28, u1_K14_29, u1_K14_30, u1_K14_31, u1_K14_32, u1_K14_33, u1_K14_34, u1_K14_35, u1_K14_36, 
       u1_K2_25, u1_K2_26, u1_K2_27, u1_K2_28, u1_K2_29, u1_K2_30, u1_K2_37, u1_K2_38, u1_K2_39, 
       u1_K2_40, u1_K2_41, u1_K2_42, u1_K3_1, u1_K3_10, u1_K3_11, u1_K3_12, u1_K3_13, u1_K3_14, 
       u1_K3_15, u1_K3_16, u1_K3_17, u1_K3_18, u1_K3_19, u1_K3_2, u1_K3_20, u1_K3_21, u1_K3_22, 
       u1_K3_23, u1_K3_24, u1_K3_3, u1_K3_4, u1_K3_5, u1_K3_6, u1_K3_7, u1_K3_8, u1_K3_9, 
       u1_K5_1, u1_K5_13, u1_K5_14, u1_K5_15, u1_K5_16, u1_K5_17, u1_K5_18, u1_K5_2, u1_K5_3, 
       u1_K5_4, u1_K5_5, u1_K5_6, u1_K7_1, u1_K7_2, u1_K7_3, u1_K7_31, u1_K7_32, u1_K7_33, 
       u1_K7_34, u1_K7_35, u1_K7_36, u1_K7_4, u1_K7_5, u1_K7_6, u1_K8_25, u1_K8_26, u1_K8_27, 
       u1_K8_28, u1_K8_29, u1_K8_30, u1_K8_31, u1_K8_32, u1_K8_33, u1_K8_34, u1_K8_35, u1_K8_36, 
       u1_K9_25, u1_K9_26, u1_K9_27, u1_K9_28, u1_K9_29, u1_K9_30, u1_out12_12, u1_out12_15, u1_out12_16, 
       u1_out12_21, u1_out12_22, u1_out12_24, u1_out12_27, u1_out12_30, u1_out12_32, u1_out12_5, u1_out12_6, u1_out12_7, 
       u1_out13_11, u1_out13_14, u1_out13_19, u1_out13_25, u1_out13_29, u1_out13_3, u1_out13_4, u1_out13_8, u1_out1_12, 
       u1_out1_14, u1_out1_22, u1_out1_25, u1_out1_3, u1_out1_32, u1_out1_7, u1_out1_8, u1_out2_1, u1_out2_10, 
       u1_out2_13, u1_out2_16, u1_out2_17, u1_out2_18, u1_out2_2, u1_out2_20, u1_out2_23, u1_out2_24, u1_out2_26, 
       u1_out2_28, u1_out2_30, u1_out2_31, u1_out2_6, u1_out2_9, u1_out4_16, u1_out4_17, u1_out4_23, u1_out4_24, 
       u1_out4_30, u1_out4_31, u1_out4_6, u1_out4_9, u1_out6_11, u1_out6_17, u1_out6_19, u1_out6_23, u1_out6_29, 
       u1_out6_31, u1_out6_4, u1_out6_9, u1_out7_11, u1_out7_14, u1_out7_19, u1_out7_25, u1_out7_29, u1_out7_3, 
       u1_out7_4, u1_out7_8, u1_out8_14, u1_out8_25, u1_out8_3, u1_out8_8, u1_out9_14, u1_out9_25, u1_out9_3, 
       u1_out9_8, u1_u12_X_13, u1_u12_X_14, u1_u12_X_15, u1_u12_X_16, u1_u12_X_17, u1_u12_X_18, u1_u12_X_37, u1_u12_X_38, 
       u1_u12_X_39, u1_u12_X_40, u1_u12_X_41, u1_u12_X_42, u1_u12_X_43, u1_u12_X_44, u1_u12_X_45, u1_u12_X_46, u1_u12_X_47, 
       u1_u12_X_48, u1_u12_u2_n100, u1_u12_u2_n101, u1_u12_u2_n102, u1_u12_u2_n103, u1_u12_u2_n104, u1_u12_u2_n105, u1_u12_u2_n106, u1_u12_u2_n107, 
       u1_u12_u2_n108, u1_u12_u2_n109, u1_u12_u2_n110, u1_u12_u2_n111, u1_u12_u2_n112, u1_u12_u2_n113, u1_u12_u2_n114, u1_u12_u2_n115, u1_u12_u2_n116, 
       u1_u12_u2_n117, u1_u12_u2_n118, u1_u12_u2_n119, u1_u12_u2_n120, u1_u12_u2_n121, u1_u12_u2_n122, u1_u12_u2_n123, u1_u12_u2_n124, u1_u12_u2_n125, 
       u1_u12_u2_n126, u1_u12_u2_n127, u1_u12_u2_n128, u1_u12_u2_n129, u1_u12_u2_n130, u1_u12_u2_n131, u1_u12_u2_n132, u1_u12_u2_n133, u1_u12_u2_n134, 
       u1_u12_u2_n135, u1_u12_u2_n136, u1_u12_u2_n137, u1_u12_u2_n138, u1_u12_u2_n139, u1_u12_u2_n140, u1_u12_u2_n141, u1_u12_u2_n142, u1_u12_u2_n143, 
       u1_u12_u2_n144, u1_u12_u2_n145, u1_u12_u2_n146, u1_u12_u2_n147, u1_u12_u2_n148, u1_u12_u2_n149, u1_u12_u2_n150, u1_u12_u2_n151, u1_u12_u2_n152, 
       u1_u12_u2_n153, u1_u12_u2_n154, u1_u12_u2_n155, u1_u12_u2_n156, u1_u12_u2_n157, u1_u12_u2_n158, u1_u12_u2_n159, u1_u12_u2_n160, u1_u12_u2_n161, 
       u1_u12_u2_n162, u1_u12_u2_n163, u1_u12_u2_n164, u1_u12_u2_n165, u1_u12_u2_n166, u1_u12_u2_n167, u1_u12_u2_n168, u1_u12_u2_n169, u1_u12_u2_n170, 
       u1_u12_u2_n171, u1_u12_u2_n172, u1_u12_u2_n173, u1_u12_u2_n174, u1_u12_u2_n175, u1_u12_u2_n176, u1_u12_u2_n177, u1_u12_u2_n178, u1_u12_u2_n179, 
       u1_u12_u2_n180, u1_u12_u2_n181, u1_u12_u2_n182, u1_u12_u2_n183, u1_u12_u2_n184, u1_u12_u2_n185, u1_u12_u2_n186, u1_u12_u2_n187, u1_u12_u2_n188, 
       u1_u12_u2_n95, u1_u12_u2_n96, u1_u12_u2_n97, u1_u12_u2_n98, u1_u12_u2_n99, u1_u12_u6_n100, u1_u12_u6_n101, u1_u12_u6_n102, u1_u12_u6_n103, 
       u1_u12_u6_n104, u1_u12_u6_n105, u1_u12_u6_n106, u1_u12_u6_n107, u1_u12_u6_n108, u1_u12_u6_n109, u1_u12_u6_n110, u1_u12_u6_n111, u1_u12_u6_n112, 
       u1_u12_u6_n113, u1_u12_u6_n114, u1_u12_u6_n115, u1_u12_u6_n116, u1_u12_u6_n117, u1_u12_u6_n118, u1_u12_u6_n119, u1_u12_u6_n120, u1_u12_u6_n121, 
       u1_u12_u6_n122, u1_u12_u6_n123, u1_u12_u6_n124, u1_u12_u6_n125, u1_u12_u6_n126, u1_u12_u6_n127, u1_u12_u6_n128, u1_u12_u6_n129, u1_u12_u6_n130, 
       u1_u12_u6_n131, u1_u12_u6_n132, u1_u12_u6_n133, u1_u12_u6_n134, u1_u12_u6_n135, u1_u12_u6_n136, u1_u12_u6_n137, u1_u12_u6_n138, u1_u12_u6_n139, 
       u1_u12_u6_n140, u1_u12_u6_n141, u1_u12_u6_n142, u1_u12_u6_n143, u1_u12_u6_n144, u1_u12_u6_n145, u1_u12_u6_n146, u1_u12_u6_n147, u1_u12_u6_n148, 
       u1_u12_u6_n149, u1_u12_u6_n150, u1_u12_u6_n151, u1_u12_u6_n152, u1_u12_u6_n153, u1_u12_u6_n154, u1_u12_u6_n155, u1_u12_u6_n156, u1_u12_u6_n157, 
       u1_u12_u6_n158, u1_u12_u6_n159, u1_u12_u6_n160, u1_u12_u6_n161, u1_u12_u6_n162, u1_u12_u6_n163, u1_u12_u6_n164, u1_u12_u6_n165, u1_u12_u6_n166, 
       u1_u12_u6_n167, u1_u12_u6_n168, u1_u12_u6_n169, u1_u12_u6_n170, u1_u12_u6_n171, u1_u12_u6_n172, u1_u12_u6_n173, u1_u12_u6_n174, u1_u12_u6_n88, 
       u1_u12_u6_n89, u1_u12_u6_n90, u1_u12_u6_n91, u1_u12_u6_n92, u1_u12_u6_n93, u1_u12_u6_n94, u1_u12_u6_n95, u1_u12_u6_n96, u1_u12_u6_n97, 
       u1_u12_u6_n98, u1_u12_u6_n99, u1_u12_u7_n100, u1_u12_u7_n101, u1_u12_u7_n102, u1_u12_u7_n103, u1_u12_u7_n104, u1_u12_u7_n105, u1_u12_u7_n106, 
       u1_u12_u7_n107, u1_u12_u7_n108, u1_u12_u7_n109, u1_u12_u7_n110, u1_u12_u7_n111, u1_u12_u7_n112, u1_u12_u7_n113, u1_u12_u7_n114, u1_u12_u7_n115, 
       u1_u12_u7_n116, u1_u12_u7_n117, u1_u12_u7_n118, u1_u12_u7_n119, u1_u12_u7_n120, u1_u12_u7_n121, u1_u12_u7_n122, u1_u12_u7_n123, u1_u12_u7_n124, 
       u1_u12_u7_n125, u1_u12_u7_n126, u1_u12_u7_n127, u1_u12_u7_n128, u1_u12_u7_n129, u1_u12_u7_n130, u1_u12_u7_n131, u1_u12_u7_n132, u1_u12_u7_n133, 
       u1_u12_u7_n134, u1_u12_u7_n135, u1_u12_u7_n136, u1_u12_u7_n137, u1_u12_u7_n138, u1_u12_u7_n139, u1_u12_u7_n140, u1_u12_u7_n141, u1_u12_u7_n142, 
       u1_u12_u7_n143, u1_u12_u7_n144, u1_u12_u7_n145, u1_u12_u7_n146, u1_u12_u7_n147, u1_u12_u7_n148, u1_u12_u7_n149, u1_u12_u7_n150, u1_u12_u7_n151, 
       u1_u12_u7_n152, u1_u12_u7_n153, u1_u12_u7_n154, u1_u12_u7_n155, u1_u12_u7_n156, u1_u12_u7_n157, u1_u12_u7_n158, u1_u12_u7_n159, u1_u12_u7_n160, 
       u1_u12_u7_n161, u1_u12_u7_n162, u1_u12_u7_n163, u1_u12_u7_n164, u1_u12_u7_n165, u1_u12_u7_n166, u1_u12_u7_n167, u1_u12_u7_n168, u1_u12_u7_n169, 
       u1_u12_u7_n170, u1_u12_u7_n171, u1_u12_u7_n172, u1_u12_u7_n173, u1_u12_u7_n174, u1_u12_u7_n175, u1_u12_u7_n176, u1_u12_u7_n177, u1_u12_u7_n178, 
       u1_u12_u7_n179, u1_u12_u7_n180, u1_u12_u7_n91, u1_u12_u7_n92, u1_u12_u7_n93, u1_u12_u7_n94, u1_u12_u7_n95, u1_u12_u7_n96, u1_u12_u7_n97, 
       u1_u12_u7_n98, u1_u12_u7_n99, u1_u13_X_25, u1_u13_X_26, u1_u13_X_27, u1_u13_X_28, u1_u13_X_29, u1_u13_X_30, u1_u13_X_31, 
       u1_u13_X_32, u1_u13_X_33, u1_u13_X_34, u1_u13_X_35, u1_u13_X_36, u1_u13_u4_n100, u1_u13_u4_n101, u1_u13_u4_n102, u1_u13_u4_n103, 
       u1_u13_u4_n104, u1_u13_u4_n105, u1_u13_u4_n106, u1_u13_u4_n107, u1_u13_u4_n108, u1_u13_u4_n109, u1_u13_u4_n110, u1_u13_u4_n111, u1_u13_u4_n112, 
       u1_u13_u4_n113, u1_u13_u4_n114, u1_u13_u4_n115, u1_u13_u4_n116, u1_u13_u4_n117, u1_u13_u4_n118, u1_u13_u4_n119, u1_u13_u4_n120, u1_u13_u4_n121, 
       u1_u13_u4_n122, u1_u13_u4_n123, u1_u13_u4_n124, u1_u13_u4_n125, u1_u13_u4_n126, u1_u13_u4_n127, u1_u13_u4_n128, u1_u13_u4_n129, u1_u13_u4_n130, 
       u1_u13_u4_n131, u1_u13_u4_n132, u1_u13_u4_n133, u1_u13_u4_n134, u1_u13_u4_n135, u1_u13_u4_n136, u1_u13_u4_n137, u1_u13_u4_n138, u1_u13_u4_n139, 
       u1_u13_u4_n140, u1_u13_u4_n141, u1_u13_u4_n142, u1_u13_u4_n143, u1_u13_u4_n144, u1_u13_u4_n145, u1_u13_u4_n146, u1_u13_u4_n147, u1_u13_u4_n148, 
       u1_u13_u4_n149, u1_u13_u4_n150, u1_u13_u4_n151, u1_u13_u4_n152, u1_u13_u4_n153, u1_u13_u4_n154, u1_u13_u4_n155, u1_u13_u4_n156, u1_u13_u4_n157, 
       u1_u13_u4_n158, u1_u13_u4_n159, u1_u13_u4_n160, u1_u13_u4_n161, u1_u13_u4_n162, u1_u13_u4_n163, u1_u13_u4_n164, u1_u13_u4_n165, u1_u13_u4_n166, 
       u1_u13_u4_n167, u1_u13_u4_n168, u1_u13_u4_n169, u1_u13_u4_n170, u1_u13_u4_n171, u1_u13_u4_n172, u1_u13_u4_n173, u1_u13_u4_n174, u1_u13_u4_n175, 
       u1_u13_u4_n176, u1_u13_u4_n177, u1_u13_u4_n178, u1_u13_u4_n179, u1_u13_u4_n180, u1_u13_u4_n181, u1_u13_u4_n182, u1_u13_u4_n183, u1_u13_u4_n184, 
       u1_u13_u4_n185, u1_u13_u4_n186, u1_u13_u4_n94, u1_u13_u4_n95, u1_u13_u4_n96, u1_u13_u4_n97, u1_u13_u4_n98, u1_u13_u4_n99, u1_u13_u5_n100, 
       u1_u13_u5_n101, u1_u13_u5_n102, u1_u13_u5_n103, u1_u13_u5_n104, u1_u13_u5_n105, u1_u13_u5_n106, u1_u13_u5_n107, u1_u13_u5_n108, u1_u13_u5_n109, 
       u1_u13_u5_n110, u1_u13_u5_n111, u1_u13_u5_n112, u1_u13_u5_n113, u1_u13_u5_n114, u1_u13_u5_n115, u1_u13_u5_n116, u1_u13_u5_n117, u1_u13_u5_n118, 
       u1_u13_u5_n119, u1_u13_u5_n120, u1_u13_u5_n121, u1_u13_u5_n122, u1_u13_u5_n123, u1_u13_u5_n124, u1_u13_u5_n125, u1_u13_u5_n126, u1_u13_u5_n127, 
       u1_u13_u5_n128, u1_u13_u5_n129, u1_u13_u5_n130, u1_u13_u5_n131, u1_u13_u5_n132, u1_u13_u5_n133, u1_u13_u5_n134, u1_u13_u5_n135, u1_u13_u5_n136, 
       u1_u13_u5_n137, u1_u13_u5_n138, u1_u13_u5_n139, u1_u13_u5_n140, u1_u13_u5_n141, u1_u13_u5_n142, u1_u13_u5_n143, u1_u13_u5_n144, u1_u13_u5_n145, 
       u1_u13_u5_n146, u1_u13_u5_n147, u1_u13_u5_n148, u1_u13_u5_n149, u1_u13_u5_n150, u1_u13_u5_n151, u1_u13_u5_n152, u1_u13_u5_n153, u1_u13_u5_n154, 
       u1_u13_u5_n155, u1_u13_u5_n156, u1_u13_u5_n157, u1_u13_u5_n158, u1_u13_u5_n159, u1_u13_u5_n160, u1_u13_u5_n161, u1_u13_u5_n162, u1_u13_u5_n163, 
       u1_u13_u5_n164, u1_u13_u5_n165, u1_u13_u5_n166, u1_u13_u5_n167, u1_u13_u5_n168, u1_u13_u5_n169, u1_u13_u5_n170, u1_u13_u5_n171, u1_u13_u5_n172, 
       u1_u13_u5_n173, u1_u13_u5_n174, u1_u13_u5_n175, u1_u13_u5_n176, u1_u13_u5_n177, u1_u13_u5_n178, u1_u13_u5_n179, u1_u13_u5_n180, u1_u13_u5_n181, 
       u1_u13_u5_n182, u1_u13_u5_n183, u1_u13_u5_n184, u1_u13_u5_n185, u1_u13_u5_n186, u1_u13_u5_n187, u1_u13_u5_n188, u1_u13_u5_n189, u1_u13_u5_n190, 
       u1_u13_u5_n191, u1_u13_u5_n192, u1_u13_u5_n193, u1_u13_u5_n194, u1_u13_u5_n195, u1_u13_u5_n196, u1_u13_u5_n99, u1_u1_X_25, u1_u1_X_26, 
       u1_u1_X_27, u1_u1_X_28, u1_u1_X_29, u1_u1_X_30, u1_u1_X_37, u1_u1_X_38, u1_u1_X_39, u1_u1_X_40, u1_u1_X_41, 
       u1_u1_X_42, u1_u1_u4_n100, u1_u1_u4_n101, u1_u1_u4_n102, u1_u1_u4_n103, u1_u1_u4_n104, u1_u1_u4_n105, u1_u1_u4_n106, u1_u1_u4_n107, 
       u1_u1_u4_n108, u1_u1_u4_n109, u1_u1_u4_n110, u1_u1_u4_n111, u1_u1_u4_n112, u1_u1_u4_n113, u1_u1_u4_n114, u1_u1_u4_n115, u1_u1_u4_n116, 
       u1_u1_u4_n117, u1_u1_u4_n118, u1_u1_u4_n119, u1_u1_u4_n120, u1_u1_u4_n121, u1_u1_u4_n122, u1_u1_u4_n123, u1_u1_u4_n124, u1_u1_u4_n125, 
       u1_u1_u4_n126, u1_u1_u4_n127, u1_u1_u4_n128, u1_u1_u4_n129, u1_u1_u4_n130, u1_u1_u4_n131, u1_u1_u4_n132, u1_u1_u4_n133, u1_u1_u4_n134, 
       u1_u1_u4_n135, u1_u1_u4_n136, u1_u1_u4_n137, u1_u1_u4_n138, u1_u1_u4_n139, u1_u1_u4_n140, u1_u1_u4_n141, u1_u1_u4_n142, u1_u1_u4_n143, 
       u1_u1_u4_n144, u1_u1_u4_n145, u1_u1_u4_n146, u1_u1_u4_n147, u1_u1_u4_n148, u1_u1_u4_n149, u1_u1_u4_n150, u1_u1_u4_n151, u1_u1_u4_n152, 
       u1_u1_u4_n153, u1_u1_u4_n154, u1_u1_u4_n155, u1_u1_u4_n156, u1_u1_u4_n157, u1_u1_u4_n158, u1_u1_u4_n159, u1_u1_u4_n160, u1_u1_u4_n161, 
       u1_u1_u4_n162, u1_u1_u4_n163, u1_u1_u4_n164, u1_u1_u4_n165, u1_u1_u4_n166, u1_u1_u4_n167, u1_u1_u4_n168, u1_u1_u4_n169, u1_u1_u4_n170, 
       u1_u1_u4_n171, u1_u1_u4_n172, u1_u1_u4_n173, u1_u1_u4_n174, u1_u1_u4_n175, u1_u1_u4_n176, u1_u1_u4_n177, u1_u1_u4_n178, u1_u1_u4_n179, 
       u1_u1_u4_n180, u1_u1_u4_n181, u1_u1_u4_n182, u1_u1_u4_n183, u1_u1_u4_n184, u1_u1_u4_n185, u1_u1_u4_n186, u1_u1_u4_n94, u1_u1_u4_n95, 
       u1_u1_u4_n96, u1_u1_u4_n97, u1_u1_u4_n98, u1_u1_u4_n99, u1_u1_u6_n100, u1_u1_u6_n101, u1_u1_u6_n102, u1_u1_u6_n103, u1_u1_u6_n104, 
       u1_u1_u6_n105, u1_u1_u6_n106, u1_u1_u6_n107, u1_u1_u6_n108, u1_u1_u6_n109, u1_u1_u6_n110, u1_u1_u6_n111, u1_u1_u6_n112, u1_u1_u6_n113, 
       u1_u1_u6_n114, u1_u1_u6_n115, u1_u1_u6_n116, u1_u1_u6_n117, u1_u1_u6_n118, u1_u1_u6_n119, u1_u1_u6_n120, u1_u1_u6_n121, u1_u1_u6_n122, 
       u1_u1_u6_n123, u1_u1_u6_n124, u1_u1_u6_n125, u1_u1_u6_n126, u1_u1_u6_n127, u1_u1_u6_n128, u1_u1_u6_n129, u1_u1_u6_n130, u1_u1_u6_n131, 
       u1_u1_u6_n132, u1_u1_u6_n133, u1_u1_u6_n134, u1_u1_u6_n135, u1_u1_u6_n136, u1_u1_u6_n137, u1_u1_u6_n138, u1_u1_u6_n139, u1_u1_u6_n140, 
       u1_u1_u6_n141, u1_u1_u6_n142, u1_u1_u6_n143, u1_u1_u6_n144, u1_u1_u6_n145, u1_u1_u6_n146, u1_u1_u6_n147, u1_u1_u6_n148, u1_u1_u6_n149, 
       u1_u1_u6_n150, u1_u1_u6_n151, u1_u1_u6_n152, u1_u1_u6_n153, u1_u1_u6_n154, u1_u1_u6_n155, u1_u1_u6_n156, u1_u1_u6_n157, u1_u1_u6_n158, 
       u1_u1_u6_n159, u1_u1_u6_n160, u1_u1_u6_n161, u1_u1_u6_n162, u1_u1_u6_n163, u1_u1_u6_n164, u1_u1_u6_n165, u1_u1_u6_n166, u1_u1_u6_n167, 
       u1_u1_u6_n168, u1_u1_u6_n169, u1_u1_u6_n170, u1_u1_u6_n171, u1_u1_u6_n172, u1_u1_u6_n173, u1_u1_u6_n174, u1_u1_u6_n88, u1_u1_u6_n89, 
       u1_u1_u6_n90, u1_u1_u6_n91, u1_u1_u6_n92, u1_u1_u6_n93, u1_u1_u6_n94, u1_u1_u6_n95, u1_u1_u6_n96, u1_u1_u6_n97, u1_u1_u6_n98, 
       u1_u1_u6_n99, u1_u2_X_1, u1_u2_X_10, u1_u2_X_11, u1_u2_X_12, u1_u2_X_13, u1_u2_X_14, u1_u2_X_15, u1_u2_X_16, 
       u1_u2_X_17, u1_u2_X_18, u1_u2_X_19, u1_u2_X_2, u1_u2_X_20, u1_u2_X_21, u1_u2_X_22, u1_u2_X_23, u1_u2_X_24, 
       u1_u2_X_3, u1_u2_X_4, u1_u2_X_5, u1_u2_X_6, u1_u2_X_7, u1_u2_X_8, u1_u2_X_9, u1_u2_u0_n100, u1_u2_u0_n101, 
       u1_u2_u0_n102, u1_u2_u0_n103, u1_u2_u0_n104, u1_u2_u0_n105, u1_u2_u0_n106, u1_u2_u0_n107, u1_u2_u0_n108, u1_u2_u0_n109, u1_u2_u0_n110, 
       u1_u2_u0_n111, u1_u2_u0_n112, u1_u2_u0_n113, u1_u2_u0_n114, u1_u2_u0_n115, u1_u2_u0_n116, u1_u2_u0_n117, u1_u2_u0_n118, u1_u2_u0_n119, 
       u1_u2_u0_n120, u1_u2_u0_n121, u1_u2_u0_n122, u1_u2_u0_n123, u1_u2_u0_n124, u1_u2_u0_n125, u1_u2_u0_n126, u1_u2_u0_n127, u1_u2_u0_n128, 
       u1_u2_u0_n129, u1_u2_u0_n130, u1_u2_u0_n131, u1_u2_u0_n132, u1_u2_u0_n133, u1_u2_u0_n134, u1_u2_u0_n135, u1_u2_u0_n136, u1_u2_u0_n137, 
       u1_u2_u0_n138, u1_u2_u0_n139, u1_u2_u0_n140, u1_u2_u0_n141, u1_u2_u0_n142, u1_u2_u0_n143, u1_u2_u0_n144, u1_u2_u0_n145, u1_u2_u0_n146, 
       u1_u2_u0_n147, u1_u2_u0_n148, u1_u2_u0_n149, u1_u2_u0_n150, u1_u2_u0_n151, u1_u2_u0_n152, u1_u2_u0_n153, u1_u2_u0_n154, u1_u2_u0_n155, 
       u1_u2_u0_n156, u1_u2_u0_n157, u1_u2_u0_n158, u1_u2_u0_n159, u1_u2_u0_n160, u1_u2_u0_n161, u1_u2_u0_n162, u1_u2_u0_n163, u1_u2_u0_n164, 
       u1_u2_u0_n165, u1_u2_u0_n166, u1_u2_u0_n167, u1_u2_u0_n168, u1_u2_u0_n169, u1_u2_u0_n170, u1_u2_u0_n171, u1_u2_u0_n172, u1_u2_u0_n173, 
       u1_u2_u0_n174, u1_u2_u0_n88, u1_u2_u0_n89, u1_u2_u0_n90, u1_u2_u0_n91, u1_u2_u0_n92, u1_u2_u0_n93, u1_u2_u0_n94, u1_u2_u0_n95, 
       u1_u2_u0_n96, u1_u2_u0_n97, u1_u2_u0_n98, u1_u2_u0_n99, u1_u2_u1_n100, u1_u2_u1_n101, u1_u2_u1_n102, u1_u2_u1_n103, u1_u2_u1_n104, 
       u1_u2_u1_n105, u1_u2_u1_n106, u1_u2_u1_n107, u1_u2_u1_n108, u1_u2_u1_n109, u1_u2_u1_n110, u1_u2_u1_n111, u1_u2_u1_n112, u1_u2_u1_n113, 
       u1_u2_u1_n114, u1_u2_u1_n115, u1_u2_u1_n116, u1_u2_u1_n117, u1_u2_u1_n118, u1_u2_u1_n119, u1_u2_u1_n120, u1_u2_u1_n121, u1_u2_u1_n122, 
       u1_u2_u1_n123, u1_u2_u1_n124, u1_u2_u1_n125, u1_u2_u1_n126, u1_u2_u1_n127, u1_u2_u1_n128, u1_u2_u1_n129, u1_u2_u1_n130, u1_u2_u1_n131, 
       u1_u2_u1_n132, u1_u2_u1_n133, u1_u2_u1_n134, u1_u2_u1_n135, u1_u2_u1_n136, u1_u2_u1_n137, u1_u2_u1_n138, u1_u2_u1_n139, u1_u2_u1_n140, 
       u1_u2_u1_n141, u1_u2_u1_n142, u1_u2_u1_n143, u1_u2_u1_n144, u1_u2_u1_n145, u1_u2_u1_n146, u1_u2_u1_n147, u1_u2_u1_n148, u1_u2_u1_n149, 
       u1_u2_u1_n150, u1_u2_u1_n151, u1_u2_u1_n152, u1_u2_u1_n153, u1_u2_u1_n154, u1_u2_u1_n155, u1_u2_u1_n156, u1_u2_u1_n157, u1_u2_u1_n158, 
       u1_u2_u1_n159, u1_u2_u1_n160, u1_u2_u1_n161, u1_u2_u1_n162, u1_u2_u1_n163, u1_u2_u1_n164, u1_u2_u1_n165, u1_u2_u1_n166, u1_u2_u1_n167, 
       u1_u2_u1_n168, u1_u2_u1_n169, u1_u2_u1_n170, u1_u2_u1_n171, u1_u2_u1_n172, u1_u2_u1_n173, u1_u2_u1_n174, u1_u2_u1_n175, u1_u2_u1_n176, 
       u1_u2_u1_n177, u1_u2_u1_n178, u1_u2_u1_n179, u1_u2_u1_n180, u1_u2_u1_n181, u1_u2_u1_n182, u1_u2_u1_n183, u1_u2_u1_n184, u1_u2_u1_n185, 
       u1_u2_u1_n186, u1_u2_u1_n187, u1_u2_u1_n188, u1_u2_u1_n95, u1_u2_u1_n96, u1_u2_u1_n97, u1_u2_u1_n98, u1_u2_u1_n99, u1_u2_u2_n100, 
       u1_u2_u2_n101, u1_u2_u2_n102, u1_u2_u2_n103, u1_u2_u2_n104, u1_u2_u2_n105, u1_u2_u2_n106, u1_u2_u2_n107, u1_u2_u2_n108, u1_u2_u2_n109, 
       u1_u2_u2_n110, u1_u2_u2_n111, u1_u2_u2_n112, u1_u2_u2_n113, u1_u2_u2_n114, u1_u2_u2_n115, u1_u2_u2_n116, u1_u2_u2_n117, u1_u2_u2_n118, 
       u1_u2_u2_n119, u1_u2_u2_n120, u1_u2_u2_n121, u1_u2_u2_n122, u1_u2_u2_n123, u1_u2_u2_n124, u1_u2_u2_n125, u1_u2_u2_n126, u1_u2_u2_n127, 
       u1_u2_u2_n128, u1_u2_u2_n129, u1_u2_u2_n130, u1_u2_u2_n131, u1_u2_u2_n132, u1_u2_u2_n133, u1_u2_u2_n134, u1_u2_u2_n135, u1_u2_u2_n136, 
       u1_u2_u2_n137, u1_u2_u2_n138, u1_u2_u2_n139, u1_u2_u2_n140, u1_u2_u2_n141, u1_u2_u2_n142, u1_u2_u2_n143, u1_u2_u2_n144, u1_u2_u2_n145, 
       u1_u2_u2_n146, u1_u2_u2_n147, u1_u2_u2_n148, u1_u2_u2_n149, u1_u2_u2_n150, u1_u2_u2_n151, u1_u2_u2_n152, u1_u2_u2_n153, u1_u2_u2_n154, 
       u1_u2_u2_n155, u1_u2_u2_n156, u1_u2_u2_n157, u1_u2_u2_n158, u1_u2_u2_n159, u1_u2_u2_n160, u1_u2_u2_n161, u1_u2_u2_n162, u1_u2_u2_n163, 
       u1_u2_u2_n164, u1_u2_u2_n165, u1_u2_u2_n166, u1_u2_u2_n167, u1_u2_u2_n168, u1_u2_u2_n169, u1_u2_u2_n170, u1_u2_u2_n171, u1_u2_u2_n172, 
       u1_u2_u2_n173, u1_u2_u2_n174, u1_u2_u2_n175, u1_u2_u2_n176, u1_u2_u2_n177, u1_u2_u2_n178, u1_u2_u2_n179, u1_u2_u2_n180, u1_u2_u2_n181, 
       u1_u2_u2_n182, u1_u2_u2_n183, u1_u2_u2_n184, u1_u2_u2_n185, u1_u2_u2_n186, u1_u2_u2_n187, u1_u2_u2_n188, u1_u2_u2_n95, u1_u2_u2_n96, 
       u1_u2_u2_n97, u1_u2_u2_n98, u1_u2_u2_n99, u1_u2_u3_n100, u1_u2_u3_n101, u1_u2_u3_n102, u1_u2_u3_n103, u1_u2_u3_n104, u1_u2_u3_n105, 
       u1_u2_u3_n106, u1_u2_u3_n107, u1_u2_u3_n108, u1_u2_u3_n109, u1_u2_u3_n110, u1_u2_u3_n111, u1_u2_u3_n112, u1_u2_u3_n113, u1_u2_u3_n114, 
       u1_u2_u3_n115, u1_u2_u3_n116, u1_u2_u3_n117, u1_u2_u3_n118, u1_u2_u3_n119, u1_u2_u3_n120, u1_u2_u3_n121, u1_u2_u3_n122, u1_u2_u3_n123, 
       u1_u2_u3_n124, u1_u2_u3_n125, u1_u2_u3_n126, u1_u2_u3_n127, u1_u2_u3_n128, u1_u2_u3_n129, u1_u2_u3_n130, u1_u2_u3_n131, u1_u2_u3_n132, 
       u1_u2_u3_n133, u1_u2_u3_n134, u1_u2_u3_n135, u1_u2_u3_n136, u1_u2_u3_n137, u1_u2_u3_n138, u1_u2_u3_n139, u1_u2_u3_n140, u1_u2_u3_n141, 
       u1_u2_u3_n142, u1_u2_u3_n143, u1_u2_u3_n144, u1_u2_u3_n145, u1_u2_u3_n146, u1_u2_u3_n147, u1_u2_u3_n148, u1_u2_u3_n149, u1_u2_u3_n150, 
       u1_u2_u3_n151, u1_u2_u3_n152, u1_u2_u3_n153, u1_u2_u3_n154, u1_u2_u3_n155, u1_u2_u3_n156, u1_u2_u3_n157, u1_u2_u3_n158, u1_u2_u3_n159, 
       u1_u2_u3_n160, u1_u2_u3_n161, u1_u2_u3_n162, u1_u2_u3_n163, u1_u2_u3_n164, u1_u2_u3_n165, u1_u2_u3_n166, u1_u2_u3_n167, u1_u2_u3_n168, 
       u1_u2_u3_n169, u1_u2_u3_n170, u1_u2_u3_n171, u1_u2_u3_n172, u1_u2_u3_n173, u1_u2_u3_n174, u1_u2_u3_n175, u1_u2_u3_n176, u1_u2_u3_n177, 
       u1_u2_u3_n178, u1_u2_u3_n179, u1_u2_u3_n180, u1_u2_u3_n181, u1_u2_u3_n182, u1_u2_u3_n183, u1_u2_u3_n184, u1_u2_u3_n185, u1_u2_u3_n186, 
       u1_u2_u3_n94, u1_u2_u3_n95, u1_u2_u3_n96, u1_u2_u3_n97, u1_u2_u3_n98, u1_u2_u3_n99, u1_u4_X_1, u1_u4_X_13, u1_u4_X_14, 
       u1_u4_X_15, u1_u4_X_16, u1_u4_X_17, u1_u4_X_18, u1_u4_X_2, u1_u4_X_3, u1_u4_X_4, u1_u4_X_5, u1_u4_X_6, 
       u1_u4_u0_n100, u1_u4_u0_n101, u1_u4_u0_n102, u1_u4_u0_n103, u1_u4_u0_n104, u1_u4_u0_n105, u1_u4_u0_n106, u1_u4_u0_n107, u1_u4_u0_n108, 
       u1_u4_u0_n109, u1_u4_u0_n110, u1_u4_u0_n111, u1_u4_u0_n112, u1_u4_u0_n113, u1_u4_u0_n114, u1_u4_u0_n115, u1_u4_u0_n116, u1_u4_u0_n117, 
       u1_u4_u0_n118, u1_u4_u0_n119, u1_u4_u0_n120, u1_u4_u0_n121, u1_u4_u0_n122, u1_u4_u0_n123, u1_u4_u0_n124, u1_u4_u0_n125, u1_u4_u0_n126, 
       u1_u4_u0_n127, u1_u4_u0_n128, u1_u4_u0_n129, u1_u4_u0_n130, u1_u4_u0_n131, u1_u4_u0_n132, u1_u4_u0_n133, u1_u4_u0_n134, u1_u4_u0_n135, 
       u1_u4_u0_n136, u1_u4_u0_n137, u1_u4_u0_n138, u1_u4_u0_n139, u1_u4_u0_n140, u1_u4_u0_n141, u1_u4_u0_n142, u1_u4_u0_n143, u1_u4_u0_n144, 
       u1_u4_u0_n145, u1_u4_u0_n146, u1_u4_u0_n147, u1_u4_u0_n148, u1_u4_u0_n149, u1_u4_u0_n150, u1_u4_u0_n151, u1_u4_u0_n152, u1_u4_u0_n153, 
       u1_u4_u0_n154, u1_u4_u0_n155, u1_u4_u0_n156, u1_u4_u0_n157, u1_u4_u0_n158, u1_u4_u0_n159, u1_u4_u0_n160, u1_u4_u0_n161, u1_u4_u0_n162, 
       u1_u4_u0_n163, u1_u4_u0_n164, u1_u4_u0_n165, u1_u4_u0_n166, u1_u4_u0_n167, u1_u4_u0_n168, u1_u4_u0_n169, u1_u4_u0_n170, u1_u4_u0_n171, 
       u1_u4_u0_n172, u1_u4_u0_n173, u1_u4_u0_n174, u1_u4_u0_n88, u1_u4_u0_n89, u1_u4_u0_n90, u1_u4_u0_n91, u1_u4_u0_n92, u1_u4_u0_n93, 
       u1_u4_u0_n94, u1_u4_u0_n95, u1_u4_u0_n96, u1_u4_u0_n97, u1_u4_u0_n98, u1_u4_u0_n99, u1_u4_u2_n100, u1_u4_u2_n101, u1_u4_u2_n102, 
       u1_u4_u2_n103, u1_u4_u2_n104, u1_u4_u2_n105, u1_u4_u2_n106, u1_u4_u2_n107, u1_u4_u2_n108, u1_u4_u2_n109, u1_u4_u2_n110, u1_u4_u2_n111, 
       u1_u4_u2_n112, u1_u4_u2_n113, u1_u4_u2_n114, u1_u4_u2_n115, u1_u4_u2_n116, u1_u4_u2_n117, u1_u4_u2_n118, u1_u4_u2_n119, u1_u4_u2_n120, 
       u1_u4_u2_n121, u1_u4_u2_n122, u1_u4_u2_n123, u1_u4_u2_n124, u1_u4_u2_n125, u1_u4_u2_n126, u1_u4_u2_n127, u1_u4_u2_n128, u1_u4_u2_n129, 
       u1_u4_u2_n130, u1_u4_u2_n131, u1_u4_u2_n132, u1_u4_u2_n133, u1_u4_u2_n134, u1_u4_u2_n135, u1_u4_u2_n136, u1_u4_u2_n137, u1_u4_u2_n138, 
       u1_u4_u2_n139, u1_u4_u2_n140, u1_u4_u2_n141, u1_u4_u2_n142, u1_u4_u2_n143, u1_u4_u2_n144, u1_u4_u2_n145, u1_u4_u2_n146, u1_u4_u2_n147, 
       u1_u4_u2_n148, u1_u4_u2_n149, u1_u4_u2_n150, u1_u4_u2_n151, u1_u4_u2_n152, u1_u4_u2_n153, u1_u4_u2_n154, u1_u4_u2_n155, u1_u4_u2_n156, 
       u1_u4_u2_n157, u1_u4_u2_n158, u1_u4_u2_n159, u1_u4_u2_n160, u1_u4_u2_n161, u1_u4_u2_n162, u1_u4_u2_n163, u1_u4_u2_n164, u1_u4_u2_n165, 
       u1_u4_u2_n166, u1_u4_u2_n167, u1_u4_u2_n168, u1_u4_u2_n169, u1_u4_u2_n170, u1_u4_u2_n171, u1_u4_u2_n172, u1_u4_u2_n173, u1_u4_u2_n174, 
       u1_u4_u2_n175, u1_u4_u2_n176, u1_u4_u2_n177, u1_u4_u2_n178, u1_u4_u2_n179, u1_u4_u2_n180, u1_u4_u2_n181, u1_u4_u2_n182, u1_u4_u2_n183, 
       u1_u4_u2_n184, u1_u4_u2_n185, u1_u4_u2_n186, u1_u4_u2_n187, u1_u4_u2_n188, u1_u4_u2_n95, u1_u4_u2_n96, u1_u4_u2_n97, u1_u4_u2_n98, 
       u1_u4_u2_n99, u1_u6_X_1, u1_u6_X_2, u1_u6_X_3, u1_u6_X_31, u1_u6_X_32, u1_u6_X_33, u1_u6_X_34, u1_u6_X_35, 
       u1_u6_X_36, u1_u6_X_4, u1_u6_X_5, u1_u6_X_6, u1_u6_u0_n100, u1_u6_u0_n101, u1_u6_u0_n102, u1_u6_u0_n103, u1_u6_u0_n104, 
       u1_u6_u0_n105, u1_u6_u0_n106, u1_u6_u0_n107, u1_u6_u0_n108, u1_u6_u0_n109, u1_u6_u0_n110, u1_u6_u0_n111, u1_u6_u0_n112, u1_u6_u0_n113, 
       u1_u6_u0_n114, u1_u6_u0_n115, u1_u6_u0_n116, u1_u6_u0_n117, u1_u6_u0_n118, u1_u6_u0_n119, u1_u6_u0_n120, u1_u6_u0_n121, u1_u6_u0_n122, 
       u1_u6_u0_n123, u1_u6_u0_n124, u1_u6_u0_n125, u1_u6_u0_n126, u1_u6_u0_n127, u1_u6_u0_n128, u1_u6_u0_n129, u1_u6_u0_n130, u1_u6_u0_n131, 
       u1_u6_u0_n132, u1_u6_u0_n133, u1_u6_u0_n134, u1_u6_u0_n135, u1_u6_u0_n136, u1_u6_u0_n137, u1_u6_u0_n138, u1_u6_u0_n139, u1_u6_u0_n140, 
       u1_u6_u0_n141, u1_u6_u0_n142, u1_u6_u0_n143, u1_u6_u0_n144, u1_u6_u0_n145, u1_u6_u0_n146, u1_u6_u0_n147, u1_u6_u0_n148, u1_u6_u0_n149, 
       u1_u6_u0_n150, u1_u6_u0_n151, u1_u6_u0_n152, u1_u6_u0_n153, u1_u6_u0_n154, u1_u6_u0_n155, u1_u6_u0_n156, u1_u6_u0_n157, u1_u6_u0_n158, 
       u1_u6_u0_n159, u1_u6_u0_n160, u1_u6_u0_n161, u1_u6_u0_n162, u1_u6_u0_n163, u1_u6_u0_n164, u1_u6_u0_n165, u1_u6_u0_n166, u1_u6_u0_n167, 
       u1_u6_u0_n168, u1_u6_u0_n169, u1_u6_u0_n170, u1_u6_u0_n171, u1_u6_u0_n172, u1_u6_u0_n173, u1_u6_u0_n174, u1_u6_u0_n88, u1_u6_u0_n89, 
       u1_u6_u0_n90, u1_u6_u0_n91, u1_u6_u0_n92, u1_u6_u0_n93, u1_u6_u0_n94, u1_u6_u0_n95, u1_u6_u0_n96, u1_u6_u0_n97, u1_u6_u0_n98, 
       u1_u6_u0_n99, u1_u6_u5_n100, u1_u6_u5_n101, u1_u6_u5_n102, u1_u6_u5_n103, u1_u6_u5_n104, u1_u6_u5_n105, u1_u6_u5_n106, u1_u6_u5_n107, 
       u1_u6_u5_n108, u1_u6_u5_n109, u1_u6_u5_n110, u1_u6_u5_n111, u1_u6_u5_n112, u1_u6_u5_n113, u1_u6_u5_n114, u1_u6_u5_n115, u1_u6_u5_n116, 
       u1_u6_u5_n117, u1_u6_u5_n118, u1_u6_u5_n119, u1_u6_u5_n120, u1_u6_u5_n121, u1_u6_u5_n122, u1_u6_u5_n123, u1_u6_u5_n124, u1_u6_u5_n125, 
       u1_u6_u5_n126, u1_u6_u5_n127, u1_u6_u5_n128, u1_u6_u5_n129, u1_u6_u5_n130, u1_u6_u5_n131, u1_u6_u5_n132, u1_u6_u5_n133, u1_u6_u5_n134, 
       u1_u6_u5_n135, u1_u6_u5_n136, u1_u6_u5_n137, u1_u6_u5_n138, u1_u6_u5_n139, u1_u6_u5_n140, u1_u6_u5_n141, u1_u6_u5_n142, u1_u6_u5_n143, 
       u1_u6_u5_n144, u1_u6_u5_n145, u1_u6_u5_n146, u1_u6_u5_n147, u1_u6_u5_n148, u1_u6_u5_n149, u1_u6_u5_n150, u1_u6_u5_n151, u1_u6_u5_n152, 
       u1_u6_u5_n153, u1_u6_u5_n154, u1_u6_u5_n155, u1_u6_u5_n156, u1_u6_u5_n157, u1_u6_u5_n158, u1_u6_u5_n159, u1_u6_u5_n160, u1_u6_u5_n161, 
       u1_u6_u5_n162, u1_u6_u5_n163, u1_u6_u5_n164, u1_u6_u5_n165, u1_u6_u5_n166, u1_u6_u5_n167, u1_u6_u5_n168, u1_u6_u5_n169, u1_u6_u5_n170, 
       u1_u6_u5_n171, u1_u6_u5_n172, u1_u6_u5_n173, u1_u6_u5_n174, u1_u6_u5_n175, u1_u6_u5_n176, u1_u6_u5_n177, u1_u6_u5_n178, u1_u6_u5_n179, 
       u1_u6_u5_n180, u1_u6_u5_n181, u1_u6_u5_n182, u1_u6_u5_n183, u1_u6_u5_n184, u1_u6_u5_n185, u1_u6_u5_n186, u1_u6_u5_n187, u1_u6_u5_n188, 
       u1_u6_u5_n189, u1_u6_u5_n190, u1_u6_u5_n191, u1_u6_u5_n192, u1_u6_u5_n193, u1_u6_u5_n194, u1_u6_u5_n195, u1_u6_u5_n196, u1_u6_u5_n99, 
       u1_u7_X_25, u1_u7_X_26, u1_u7_X_27, u1_u7_X_28, u1_u7_X_29, u1_u7_X_30, u1_u7_X_31, u1_u7_X_32, u1_u7_X_33, 
       u1_u7_X_34, u1_u7_X_35, u1_u7_X_36, u1_u7_u4_n100, u1_u7_u4_n101, u1_u7_u4_n102, u1_u7_u4_n103, u1_u7_u4_n104, u1_u7_u4_n105, 
       u1_u7_u4_n106, u1_u7_u4_n107, u1_u7_u4_n108, u1_u7_u4_n109, u1_u7_u4_n110, u1_u7_u4_n111, u1_u7_u4_n112, u1_u7_u4_n113, u1_u7_u4_n114, 
       u1_u7_u4_n115, u1_u7_u4_n116, u1_u7_u4_n117, u1_u7_u4_n118, u1_u7_u4_n119, u1_u7_u4_n120, u1_u7_u4_n121, u1_u7_u4_n122, u1_u7_u4_n123, 
       u1_u7_u4_n124, u1_u7_u4_n125, u1_u7_u4_n126, u1_u7_u4_n127, u1_u7_u4_n128, u1_u7_u4_n129, u1_u7_u4_n130, u1_u7_u4_n131, u1_u7_u4_n132, 
       u1_u7_u4_n133, u1_u7_u4_n134, u1_u7_u4_n135, u1_u7_u4_n136, u1_u7_u4_n137, u1_u7_u4_n138, u1_u7_u4_n139, u1_u7_u4_n140, u1_u7_u4_n141, 
       u1_u7_u4_n142, u1_u7_u4_n143, u1_u7_u4_n144, u1_u7_u4_n145, u1_u7_u4_n146, u1_u7_u4_n147, u1_u7_u4_n148, u1_u7_u4_n149, u1_u7_u4_n150, 
       u1_u7_u4_n151, u1_u7_u4_n152, u1_u7_u4_n153, u1_u7_u4_n154, u1_u7_u4_n155, u1_u7_u4_n156, u1_u7_u4_n157, u1_u7_u4_n158, u1_u7_u4_n159, 
       u1_u7_u4_n160, u1_u7_u4_n161, u1_u7_u4_n162, u1_u7_u4_n163, u1_u7_u4_n164, u1_u7_u4_n165, u1_u7_u4_n166, u1_u7_u4_n167, u1_u7_u4_n168, 
       u1_u7_u4_n169, u1_u7_u4_n170, u1_u7_u4_n171, u1_u7_u4_n172, u1_u7_u4_n173, u1_u7_u4_n174, u1_u7_u4_n175, u1_u7_u4_n176, u1_u7_u4_n177, 
       u1_u7_u4_n178, u1_u7_u4_n179, u1_u7_u4_n180, u1_u7_u4_n181, u1_u7_u4_n182, u1_u7_u4_n183, u1_u7_u4_n184, u1_u7_u4_n185, u1_u7_u4_n186, 
       u1_u7_u4_n94, u1_u7_u4_n95, u1_u7_u4_n96, u1_u7_u4_n97, u1_u7_u4_n98, u1_u7_u4_n99, u1_u7_u5_n100, u1_u7_u5_n101, u1_u7_u5_n102, 
       u1_u7_u5_n103, u1_u7_u5_n104, u1_u7_u5_n105, u1_u7_u5_n106, u1_u7_u5_n107, u1_u7_u5_n108, u1_u7_u5_n109, u1_u7_u5_n110, u1_u7_u5_n111, 
       u1_u7_u5_n112, u1_u7_u5_n113, u1_u7_u5_n114, u1_u7_u5_n115, u1_u7_u5_n116, u1_u7_u5_n117, u1_u7_u5_n118, u1_u7_u5_n119, u1_u7_u5_n120, 
       u1_u7_u5_n121, u1_u7_u5_n122, u1_u7_u5_n123, u1_u7_u5_n124, u1_u7_u5_n125, u1_u7_u5_n126, u1_u7_u5_n127, u1_u7_u5_n128, u1_u7_u5_n129, 
       u1_u7_u5_n130, u1_u7_u5_n131, u1_u7_u5_n132, u1_u7_u5_n133, u1_u7_u5_n134, u1_u7_u5_n135, u1_u7_u5_n136, u1_u7_u5_n137, u1_u7_u5_n138, 
       u1_u7_u5_n139, u1_u7_u5_n140, u1_u7_u5_n141, u1_u7_u5_n142, u1_u7_u5_n143, u1_u7_u5_n144, u1_u7_u5_n145, u1_u7_u5_n146, u1_u7_u5_n147, 
       u1_u7_u5_n148, u1_u7_u5_n149, u1_u7_u5_n150, u1_u7_u5_n151, u1_u7_u5_n152, u1_u7_u5_n153, u1_u7_u5_n154, u1_u7_u5_n155, u1_u7_u5_n156, 
       u1_u7_u5_n157, u1_u7_u5_n158, u1_u7_u5_n159, u1_u7_u5_n160, u1_u7_u5_n161, u1_u7_u5_n162, u1_u7_u5_n163, u1_u7_u5_n164, u1_u7_u5_n165, 
       u1_u7_u5_n166, u1_u7_u5_n167, u1_u7_u5_n168, u1_u7_u5_n169, u1_u7_u5_n170, u1_u7_u5_n171, u1_u7_u5_n172, u1_u7_u5_n173, u1_u7_u5_n174, 
       u1_u7_u5_n175, u1_u7_u5_n176, u1_u7_u5_n177, u1_u7_u5_n178, u1_u7_u5_n179, u1_u7_u5_n180, u1_u7_u5_n181, u1_u7_u5_n182, u1_u7_u5_n183, 
       u1_u7_u5_n184, u1_u7_u5_n185, u1_u7_u5_n186, u1_u7_u5_n187, u1_u7_u5_n188, u1_u7_u5_n189, u1_u7_u5_n190, u1_u7_u5_n191, u1_u7_u5_n192, 
       u1_u7_u5_n193, u1_u7_u5_n194, u1_u7_u5_n195, u1_u7_u5_n196, u1_u7_u5_n99, u1_u8_X_25, u1_u8_X_26, u1_u8_X_27, u1_u8_X_28, 
       u1_u8_X_29, u1_u8_X_30, u1_u8_u4_n100, u1_u8_u4_n101, u1_u8_u4_n102, u1_u8_u4_n103, u1_u8_u4_n104, u1_u8_u4_n105, u1_u8_u4_n106, 
       u1_u8_u4_n107, u1_u8_u4_n108, u1_u8_u4_n109, u1_u8_u4_n110, u1_u8_u4_n111, u1_u8_u4_n112, u1_u8_u4_n113, u1_u8_u4_n114, u1_u8_u4_n115, 
       u1_u8_u4_n116, u1_u8_u4_n117, u1_u8_u4_n118, u1_u8_u4_n119, u1_u8_u4_n120, u1_u8_u4_n121, u1_u8_u4_n122, u1_u8_u4_n123, u1_u8_u4_n124, 
       u1_u8_u4_n125, u1_u8_u4_n126, u1_u8_u4_n127, u1_u8_u4_n128, u1_u8_u4_n129, u1_u8_u4_n130, u1_u8_u4_n131, u1_u8_u4_n132, u1_u8_u4_n133, 
       u1_u8_u4_n134, u1_u8_u4_n135, u1_u8_u4_n136, u1_u8_u4_n137, u1_u8_u4_n138, u1_u8_u4_n139, u1_u8_u4_n140, u1_u8_u4_n141, u1_u8_u4_n142, 
       u1_u8_u4_n143, u1_u8_u4_n144, u1_u8_u4_n145, u1_u8_u4_n146, u1_u8_u4_n147, u1_u8_u4_n148, u1_u8_u4_n149, u1_u8_u4_n150, u1_u8_u4_n151, 
       u1_u8_u4_n152, u1_u8_u4_n153, u1_u8_u4_n154, u1_u8_u4_n155, u1_u8_u4_n156, u1_u8_u4_n157, u1_u8_u4_n158, u1_u8_u4_n159, u1_u8_u4_n160, 
       u1_u8_u4_n161, u1_u8_u4_n162, u1_u8_u4_n163, u1_u8_u4_n164, u1_u8_u4_n165, u1_u8_u4_n166, u1_u8_u4_n167, u1_u8_u4_n168, u1_u8_u4_n169, 
       u1_u8_u4_n170, u1_u8_u4_n171, u1_u8_u4_n172, u1_u8_u4_n173, u1_u8_u4_n174, u1_u8_u4_n175, u1_u8_u4_n176, u1_u8_u4_n177, u1_u8_u4_n178, 
       u1_u8_u4_n179, u1_u8_u4_n180, u1_u8_u4_n181, u1_u8_u4_n182, u1_u8_u4_n183, u1_u8_u4_n184, u1_u8_u4_n185, u1_u8_u4_n186, u1_u8_u4_n94, 
       u1_u8_u4_n95, u1_u8_u4_n96, u1_u8_u4_n97, u1_u8_u4_n98, u1_u8_u4_n99, u1_u9_X_25, u1_u9_X_26, u1_u9_X_27, u1_u9_X_28, 
       u1_u9_X_29, u1_u9_X_30, u1_u9_u4_n100, u1_u9_u4_n101, u1_u9_u4_n102, u1_u9_u4_n103, u1_u9_u4_n104, u1_u9_u4_n105, u1_u9_u4_n106, 
       u1_u9_u4_n107, u1_u9_u4_n108, u1_u9_u4_n109, u1_u9_u4_n110, u1_u9_u4_n111, u1_u9_u4_n112, u1_u9_u4_n113, u1_u9_u4_n114, u1_u9_u4_n115, 
       u1_u9_u4_n116, u1_u9_u4_n117, u1_u9_u4_n118, u1_u9_u4_n119, u1_u9_u4_n120, u1_u9_u4_n121, u1_u9_u4_n122, u1_u9_u4_n123, u1_u9_u4_n124, 
       u1_u9_u4_n125, u1_u9_u4_n126, u1_u9_u4_n127, u1_u9_u4_n128, u1_u9_u4_n129, u1_u9_u4_n130, u1_u9_u4_n131, u1_u9_u4_n132, u1_u9_u4_n133, 
       u1_u9_u4_n134, u1_u9_u4_n135, u1_u9_u4_n136, u1_u9_u4_n137, u1_u9_u4_n138, u1_u9_u4_n139, u1_u9_u4_n140, u1_u9_u4_n141, u1_u9_u4_n142, 
       u1_u9_u4_n143, u1_u9_u4_n144, u1_u9_u4_n145, u1_u9_u4_n146, u1_u9_u4_n147, u1_u9_u4_n148, u1_u9_u4_n149, u1_u9_u4_n150, u1_u9_u4_n151, 
       u1_u9_u4_n152, u1_u9_u4_n153, u1_u9_u4_n154, u1_u9_u4_n155, u1_u9_u4_n156, u1_u9_u4_n157, u1_u9_u4_n158, u1_u9_u4_n159, u1_u9_u4_n160, 
       u1_u9_u4_n161, u1_u9_u4_n162, u1_u9_u4_n163, u1_u9_u4_n164, u1_u9_u4_n165, u1_u9_u4_n166, u1_u9_u4_n167, u1_u9_u4_n168, u1_u9_u4_n169, 
       u1_u9_u4_n170, u1_u9_u4_n171, u1_u9_u4_n172, u1_u9_u4_n173, u1_u9_u4_n174, u1_u9_u4_n175, u1_u9_u4_n176, u1_u9_u4_n177, u1_u9_u4_n178, 
       u1_u9_u4_n179, u1_u9_u4_n180, u1_u9_u4_n181, u1_u9_u4_n182, u1_u9_u4_n183, u1_u9_u4_n184, u1_u9_u4_n185, u1_u9_u4_n186, u1_u9_u4_n94, 
       u1_u9_u4_n95, u1_u9_u4_n96, u1_u9_u4_n97, u1_u9_u4_n98, u1_u9_u4_n99, u1_uk_n1026, u1_uk_n1027, u1_uk_n1028, u1_uk_n1031, 
       u1_uk_n1036, u1_uk_n1037, u1_uk_n1038, u1_uk_n1043, u1_uk_n1048, u1_uk_n1049, u1_uk_n1072, u1_uk_n1085, u1_uk_n1086, 
       u1_uk_n1108, u1_uk_n1116, u1_uk_n1117, u1_uk_n1118, u1_uk_n1119, u1_uk_n1120, u1_uk_n1121, u1_uk_n1125, u1_uk_n1133, 
       u1_uk_n1134, u1_uk_n1136, u1_uk_n1137, u1_uk_n1158, u1_uk_n1159, u1_uk_n1161, u1_uk_n335, u1_uk_n677, u1_uk_n678, 
       u1_uk_n681, u1_uk_n682, u1_uk_n946, u1_uk_n947, u1_uk_n953, u1_uk_n954, u1_uk_n955, u1_uk_n956, u2_K16_43, 
       u2_K16_45, u2_K16_46, u2_K16_48, u2_K7_19, u2_K7_20, u2_K7_21, u2_K7_22, u2_K7_23, u2_K7_24, 
       u2_out15_15, u2_out15_21, u2_out15_27, u2_out15_5, u2_out6_1, u2_out6_10, u2_out6_20, u2_out6_26, u2_u15_X_43, 
       u2_u15_X_44, u2_u15_X_45, u2_u15_X_46, u2_u15_X_47, u2_u15_X_48, u2_u15_u7_n100, u2_u15_u7_n101, u2_u15_u7_n102, u2_u15_u7_n103, 
       u2_u15_u7_n104, u2_u15_u7_n105, u2_u15_u7_n106, u2_u15_u7_n107, u2_u15_u7_n108, u2_u15_u7_n109, u2_u15_u7_n110, u2_u15_u7_n111, u2_u15_u7_n112, 
       u2_u15_u7_n113, u2_u15_u7_n114, u2_u15_u7_n115, u2_u15_u7_n116, u2_u15_u7_n117, u2_u15_u7_n118, u2_u15_u7_n119, u2_u15_u7_n120, u2_u15_u7_n121, 
       u2_u15_u7_n122, u2_u15_u7_n123, u2_u15_u7_n124, u2_u15_u7_n125, u2_u15_u7_n126, u2_u15_u7_n127, u2_u15_u7_n128, u2_u15_u7_n129, u2_u15_u7_n130, 
       u2_u15_u7_n131, u2_u15_u7_n132, u2_u15_u7_n133, u2_u15_u7_n134, u2_u15_u7_n135, u2_u15_u7_n136, u2_u15_u7_n137, u2_u15_u7_n138, u2_u15_u7_n139, 
       u2_u15_u7_n140, u2_u15_u7_n141, u2_u15_u7_n142, u2_u15_u7_n143, u2_u15_u7_n144, u2_u15_u7_n145, u2_u15_u7_n146, u2_u15_u7_n147, u2_u15_u7_n148, 
       u2_u15_u7_n149, u2_u15_u7_n150, u2_u15_u7_n151, u2_u15_u7_n152, u2_u15_u7_n153, u2_u15_u7_n154, u2_u15_u7_n155, u2_u15_u7_n156, u2_u15_u7_n157, 
       u2_u15_u7_n158, u2_u15_u7_n159, u2_u15_u7_n160, u2_u15_u7_n161, u2_u15_u7_n162, u2_u15_u7_n163, u2_u15_u7_n164, u2_u15_u7_n165, u2_u15_u7_n166, 
       u2_u15_u7_n167, u2_u15_u7_n168, u2_u15_u7_n169, u2_u15_u7_n170, u2_u15_u7_n171, u2_u15_u7_n172, u2_u15_u7_n173, u2_u15_u7_n174, u2_u15_u7_n175, 
       u2_u15_u7_n176, u2_u15_u7_n177, u2_u15_u7_n178, u2_u15_u7_n179, u2_u15_u7_n180, u2_u15_u7_n91, u2_u15_u7_n92, u2_u15_u7_n93, u2_u15_u7_n94, 
       u2_u15_u7_n95, u2_u15_u7_n96, u2_u15_u7_n97, u2_u15_u7_n98, u2_u15_u7_n99, u2_u6_X_19, u2_u6_X_20, u2_u6_X_21, u2_u6_X_22, 
       u2_u6_X_23, u2_u6_X_24, u2_u6_u3_n100, u2_u6_u3_n101, u2_u6_u3_n102, u2_u6_u3_n103, u2_u6_u3_n104, u2_u6_u3_n105, u2_u6_u3_n106, 
       u2_u6_u3_n107, u2_u6_u3_n108, u2_u6_u3_n109, u2_u6_u3_n110, u2_u6_u3_n111, u2_u6_u3_n112, u2_u6_u3_n113, u2_u6_u3_n114, u2_u6_u3_n115, 
       u2_u6_u3_n116, u2_u6_u3_n117, u2_u6_u3_n118, u2_u6_u3_n119, u2_u6_u3_n120, u2_u6_u3_n121, u2_u6_u3_n122, u2_u6_u3_n123, u2_u6_u3_n124, 
       u2_u6_u3_n125, u2_u6_u3_n126, u2_u6_u3_n127, u2_u6_u3_n128, u2_u6_u3_n129, u2_u6_u3_n130, u2_u6_u3_n131, u2_u6_u3_n132, u2_u6_u3_n133, 
       u2_u6_u3_n134, u2_u6_u3_n135, u2_u6_u3_n136, u2_u6_u3_n137, u2_u6_u3_n138, u2_u6_u3_n139, u2_u6_u3_n140, u2_u6_u3_n141, u2_u6_u3_n142, 
       u2_u6_u3_n143, u2_u6_u3_n144, u2_u6_u3_n145, u2_u6_u3_n146, u2_u6_u3_n147, u2_u6_u3_n148, u2_u6_u3_n149, u2_u6_u3_n150, u2_u6_u3_n151, 
       u2_u6_u3_n152, u2_u6_u3_n153, u2_u6_u3_n154, u2_u6_u3_n155, u2_u6_u3_n156, u2_u6_u3_n157, u2_u6_u3_n158, u2_u6_u3_n159, u2_u6_u3_n160, 
       u2_u6_u3_n161, u2_u6_u3_n162, u2_u6_u3_n163, u2_u6_u3_n164, u2_u6_u3_n165, u2_u6_u3_n166, u2_u6_u3_n167, u2_u6_u3_n168, u2_u6_u3_n169, 
       u2_u6_u3_n170, u2_u6_u3_n171, u2_u6_u3_n172, u2_u6_u3_n173, u2_u6_u3_n174, u2_u6_u3_n175, u2_u6_u3_n176, u2_u6_u3_n177, u2_u6_u3_n178, 
       u2_u6_u3_n179, u2_u6_u3_n180, u2_u6_u3_n181, u2_u6_u3_n182, u2_u6_u3_n183, u2_u6_u3_n184, u2_u6_u3_n185, u2_u6_u3_n186, u2_u6_u3_n94, 
       u2_u6_u3_n95, u2_u6_u3_n96, u2_u6_u3_n97, u2_u6_u3_n98, u2_u6_u3_n99, u2_uk_n1080, u2_uk_n1083,  u2_uk_n963;
  XOR2_X1 u1_U102 (.B( u1_L12_25 ) , .Z( u1_N440 ) , .A( u1_out13_25 ) );
  XOR2_X1 u1_U109 (.B( u1_L12_19 ) , .Z( u1_N434 ) , .A( u1_out13_19 ) );
  XOR2_X1 u1_U11 (.B( u1_L1_28 ) , .Z( u1_N91 ) , .A( u1_out2_28 ) );
  XOR2_X1 u1_U114 (.B( u1_L0_12 ) , .Z( u1_N43 ) , .A( u1_out1_12 ) );
  XOR2_X1 u1_U115 (.B( u1_L12_14 ) , .Z( u1_N429 ) , .A( u1_out13_14 ) );
  XOR2_X1 u1_U118 (.B( u1_L12_11 ) , .Z( u1_N426 ) , .A( u1_out13_11 ) );
  XOR2_X1 u1_U121 (.B( u1_L12_8 ) , .Z( u1_N423 ) , .A( u1_out13_8 ) );
  XOR2_X1 u1_U126 (.B( u1_L12_4 ) , .Z( u1_N419 ) , .A( u1_out13_4 ) );
  XOR2_X1 u1_U127 (.B( u1_L12_3 ) , .Z( u1_N418 ) , .A( u1_out13_3 ) );
  XOR2_X1 u1_U130 (.B( u1_L11_32 ) , .Z( u1_N415 ) , .A( u1_out12_32 ) );
  XOR2_X1 u1_U132 (.B( u1_L11_30 ) , .Z( u1_N413 ) , .A( u1_out12_30 ) );
  XOR2_X1 u1_U135 (.B( u1_L11_27 ) , .Z( u1_N410 ) , .A( u1_out12_27 ) );
  XOR2_X1 u1_U139 (.B( u1_L11_24 ) , .Z( u1_N407 ) , .A( u1_out12_24 ) );
  XOR2_X1 u1_U14 (.B( u1_L1_26 ) , .Z( u1_N89 ) , .A( u1_out2_26 ) );
  XOR2_X1 u1_U141 (.B( u1_L11_22 ) , .Z( u1_N405 ) , .A( u1_out12_22 ) );
  XOR2_X1 u1_U142 (.B( u1_L11_21 ) , .Z( u1_N404 ) , .A( u1_out12_21 ) );
  XOR2_X1 u1_U149 (.B( u1_L11_16 ) , .Z( u1_N399 ) , .A( u1_out12_16 ) );
  XOR2_X1 u1_U150 (.B( u1_L11_15 ) , .Z( u1_N398 ) , .A( u1_out12_15 ) );
  XOR2_X1 u1_U153 (.B( u1_L11_12 ) , .Z( u1_N395 ) , .A( u1_out12_12 ) );
  XOR2_X1 u1_U158 (.B( u1_L11_7 ) , .Z( u1_N390 ) , .A( u1_out12_7 ) );
  XOR2_X1 u1_U159 (.B( u1_L0_8 ) , .Z( u1_N39 ) , .A( u1_out1_8 ) );
  XOR2_X1 u1_U16 (.B( u1_L1_24 ) , .Z( u1_N87 ) , .A( u1_out2_24 ) );
  XOR2_X1 u1_U160 (.B( u1_L11_6 ) , .Z( u1_N389 ) , .A( u1_out12_6 ) );
  XOR2_X1 u1_U161 (.B( u1_L11_5 ) , .Z( u1_N388 ) , .A( u1_out12_5 ) );
  XOR2_X1 u1_U17 (.B( u1_L1_23 ) , .Z( u1_N86 ) , .A( u1_out2_23 ) );
  XOR2_X1 u1_U170 (.B( u1_L0_7 ) , .Z( u1_N38 ) , .A( u1_out1_7 ) );
  XOR2_X1 u1_U20 (.B( u1_L1_20 ) , .Z( u1_N83 ) , .A( u1_out2_20 ) );
  XOR2_X1 u1_U214 (.B( u1_L0_3 ) , .Z( u1_N34 ) , .A( u1_out1_3 ) );
  XOR2_X1 u1_U22 (.B( u1_L1_18 ) , .Z( u1_N81 ) , .A( u1_out2_18 ) );
  XOR2_X1 u1_U23 (.B( u1_L1_17 ) , .Z( u1_N80 ) , .A( u1_out2_17 ) );
  XOR2_X1 u1_U244 (.B( u1_L8_25 ) , .Z( u1_N312 ) , .A( u1_out9_25 ) );
  XOR2_X1 u1_U25 (.B( u1_L1_16 ) , .Z( u1_N79 ) , .A( u1_out2_16 ) );
  XOR2_X1 u1_U256 (.B( u1_L8_14 ) , .Z( u1_N301 ) , .A( u1_out9_14 ) );
  XOR2_X1 u1_U264 (.B( u1_L8_8 ) , .Z( u1_N295 ) , .A( u1_out9_8 ) );
  XOR2_X1 u1_U269 (.B( u1_L8_3 ) , .Z( u1_N290 ) , .A( u1_out9_3 ) );
  XOR2_X1 u1_U28 (.B( u1_L1_13 ) , .Z( u1_N76 ) , .A( u1_out2_13 ) );
  XOR2_X1 u1_U280 (.B( u1_L7_25 ) , .Z( u1_N280 ) , .A( u1_out8_25 ) );
  XOR2_X1 u1_U293 (.B( u1_L7_14 ) , .Z( u1_N269 ) , .A( u1_out8_14 ) );
  XOR2_X1 u1_U299 (.B( u1_L7_8 ) , .Z( u1_N263 ) , .A( u1_out8_8 ) );
  XOR2_X1 u1_U305 (.B( u1_L7_3 ) , .Z( u1_N258 ) , .A( u1_out8_3 ) );
  XOR2_X1 u1_U31 (.B( u1_L1_10 ) , .Z( u1_N73 ) , .A( u1_out2_10 ) );
  XOR2_X1 u1_U311 (.B( u1_L6_29 ) , .Z( u1_N252 ) , .A( u1_out7_29 ) );
  XOR2_X1 u1_U316 (.B( u1_L6_25 ) , .Z( u1_N248 ) , .A( u1_out7_25 ) );
  XOR2_X1 u1_U32 (.B( u1_L1_9 ) , .Z( u1_N72 ) , .A( u1_out2_9 ) );
  XOR2_X1 u1_U322 (.B( u1_L6_19 ) , .Z( u1_N242 ) , .A( u1_out7_19 ) );
  XOR2_X1 u1_U328 (.B( u1_L6_14 ) , .Z( u1_N237 ) , .A( u1_out7_14 ) );
  XOR2_X1 u1_U331 (.B( u1_L6_11 ) , .Z( u1_N234 ) , .A( u1_out7_11 ) );
  XOR2_X1 u1_U334 (.B( u1_L6_8 ) , .Z( u1_N231 ) , .A( u1_out7_8 ) );
  XOR2_X1 u1_U339 (.B( u1_L6_4 ) , .Z( u1_N227 ) , .A( u1_out7_4 ) );
  XOR2_X1 u1_U340 (.B( u1_L6_3 ) , .Z( u1_N226 ) , .A( u1_out7_3 ) );
  XOR2_X1 u1_U344 (.B( u1_L5_31 ) , .Z( u1_N222 ) , .A( u1_out6_31 ) );
  XOR2_X1 u1_U346 (.B( u1_L5_29 ) , .Z( u1_N220 ) , .A( u1_out6_29 ) );
  XOR2_X1 u1_U353 (.B( u1_L5_23 ) , .Z( u1_N214 ) , .A( u1_out6_23 ) );
  XOR2_X1 u1_U357 (.B( u1_L5_19 ) , .Z( u1_N210 ) , .A( u1_out6_19 ) );
  XOR2_X1 u1_U36 (.B( u1_L1_6 ) , .Z( u1_N69 ) , .A( u1_out2_6 ) );
  XOR2_X1 u1_U360 (.B( u1_L5_17 ) , .Z( u1_N208 ) , .A( u1_out6_17 ) );
  XOR2_X1 u1_U366 (.B( u1_L5_11 ) , .Z( u1_N202 ) , .A( u1_out6_11 ) );
  XOR2_X1 u1_U368 (.B( u1_L5_9 ) , .Z( u1_N200 ) , .A( u1_out6_9 ) );
  XOR2_X1 u1_U375 (.B( u1_L5_4 ) , .Z( u1_N195 ) , .A( u1_out6_4 ) );
  XOR2_X1 u1_U40 (.B( u1_L1_2 ) , .Z( u1_N65 ) , .A( u1_out2_2 ) );
  XOR2_X1 u1_U41 (.B( u1_L1_1 ) , .Z( u1_N64 ) , .A( u1_out2_1 ) );
  XOR2_X1 u1_U416 (.B( u1_L3_31 ) , .Z( u1_N158 ) , .A( u1_out4_31 ) );
  XOR2_X1 u1_U417 (.B( u1_L3_30 ) , .Z( u1_N157 ) , .A( u1_out4_30 ) );
  XOR2_X1 u1_U42 (.B( u1_L0_32 ) , .Z( u1_N63 ) , .A( u1_out1_32 ) );
  XOR2_X1 u1_U423 (.B( u1_L3_24 ) , .Z( u1_N151 ) , .A( u1_out4_24 ) );
  XOR2_X1 u1_U424 (.B( u1_L3_23 ) , .Z( u1_N150 ) , .A( u1_out4_23 ) );
  XOR2_X1 u1_U431 (.B( u1_L3_17 ) , .Z( u1_N144 ) , .A( u1_out4_17 ) );
  XOR2_X1 u1_U432 (.B( u1_L3_16 ) , .Z( u1_N143 ) , .A( u1_out4_16 ) );
  XOR2_X1 u1_U440 (.B( u1_L3_9 ) , .Z( u1_N136 ) , .A( u1_out4_9 ) );
  XOR2_X1 u1_U443 (.B( u1_L3_6 ) , .Z( u1_N133 ) , .A( u1_out4_6 ) );
  XOR2_X1 u1_U50 (.B( u1_L0_25 ) , .Z( u1_N56 ) , .A( u1_out1_25 ) );
  XOR2_X1 u1_U53 (.B( u1_L0_22 ) , .Z( u1_N53 ) , .A( u1_out1_22 ) );
  XOR2_X1 u1_U8 (.B( u1_L1_31 ) , .Z( u1_N94 ) , .A( u1_out2_31 ) );
  XOR2_X1 u1_U9 (.B( u1_L1_30 ) , .Z( u1_N93 ) , .A( u1_out2_30 ) );
  XOR2_X1 u1_U92 (.B( u1_L0_14 ) , .Z( u1_N45 ) , .A( u1_out1_14 ) );
  XOR2_X1 u1_U98 (.B( u1_L12_29 ) , .Z( u1_N444 ) , .A( u1_out13_29 ) );
  XOR2_X1 u1_u12_U10 (.B( u1_K13_45 ) , .A( u1_R11_30 ) , .Z( u1_u12_X_45 ) );
  XOR2_X1 u1_u12_U11 (.B( u1_K13_44 ) , .A( u1_R11_29 ) , .Z( u1_u12_X_44 ) );
  XOR2_X1 u1_u12_U12 (.B( u1_K13_43 ) , .A( u1_R11_28 ) , .Z( u1_u12_X_43 ) );
  XOR2_X1 u1_u12_U13 (.B( u1_K13_42 ) , .A( u1_R11_29 ) , .Z( u1_u12_X_42 ) );
  XOR2_X1 u1_u12_U14 (.B( u1_K13_41 ) , .A( u1_R11_28 ) , .Z( u1_u12_X_41 ) );
  XOR2_X1 u1_u12_U15 (.B( u1_K13_40 ) , .A( u1_R11_27 ) , .Z( u1_u12_X_40 ) );
  XOR2_X1 u1_u12_U17 (.B( u1_K13_39 ) , .A( u1_R11_26 ) , .Z( u1_u12_X_39 ) );
  XOR2_X1 u1_u12_U18 (.B( u1_K13_38 ) , .A( u1_R11_25 ) , .Z( u1_u12_X_38 ) );
  XOR2_X1 u1_u12_U19 (.B( u1_K13_37 ) , .A( u1_R11_24 ) , .Z( u1_u12_X_37 ) );
  XOR2_X1 u1_u12_U40 (.B( u1_K13_18 ) , .A( u1_R11_13 ) , .Z( u1_u12_X_18 ) );
  XOR2_X1 u1_u12_U41 (.B( u1_K13_17 ) , .A( u1_R11_12 ) , .Z( u1_u12_X_17 ) );
  XOR2_X1 u1_u12_U42 (.B( u1_K13_16 ) , .A( u1_R11_11 ) , .Z( u1_u12_X_16 ) );
  XOR2_X1 u1_u12_U43 (.B( u1_K13_15 ) , .A( u1_R11_10 ) , .Z( u1_u12_X_15 ) );
  XOR2_X1 u1_u12_U44 (.B( u1_K13_14 ) , .A( u1_R11_9 ) , .Z( u1_u12_X_14 ) );
  XOR2_X1 u1_u12_U45 (.B( u1_K13_13 ) , .A( u1_R11_8 ) , .Z( u1_u12_X_13 ) );
  XOR2_X1 u1_u12_U7 (.B( u1_K13_48 ) , .A( u1_R11_1 ) , .Z( u1_u12_X_48 ) );
  XOR2_X1 u1_u12_U8 (.B( u1_K13_47 ) , .A( u1_R11_32 ) , .Z( u1_u12_X_47 ) );
  XOR2_X1 u1_u12_U9 (.B( u1_K13_46 ) , .A( u1_R11_31 ) , .Z( u1_u12_X_46 ) );
  OAI22_X1 u1_u12_u2_U10 (.B1( u1_u12_u2_n151 ) , .A2( u1_u12_u2_n152 ) , .A1( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n160 ) , .B2( u1_u12_u2_n168 ) );
  NAND3_X1 u1_u12_u2_U100 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n104 ) , .A3( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n98 ) );
  NOR3_X1 u1_u12_u2_U11 (.A1( u1_u12_u2_n150 ) , .ZN( u1_u12_u2_n151 ) , .A3( u1_u12_u2_n175 ) , .A2( u1_u12_u2_n188 ) );
  AOI21_X1 u1_u12_u2_U12 (.B2( u1_u12_u2_n123 ) , .ZN( u1_u12_u2_n125 ) , .A( u1_u12_u2_n171 ) , .B1( u1_u12_u2_n184 ) );
  INV_X1 u1_u12_u2_U13 (.A( u1_u12_u2_n150 ) , .ZN( u1_u12_u2_n184 ) );
  AOI21_X1 u1_u12_u2_U14 (.ZN( u1_u12_u2_n144 ) , .B2( u1_u12_u2_n155 ) , .A( u1_u12_u2_n172 ) , .B1( u1_u12_u2_n185 ) );
  AOI21_X1 u1_u12_u2_U15 (.B2( u1_u12_u2_n143 ) , .ZN( u1_u12_u2_n145 ) , .B1( u1_u12_u2_n152 ) , .A( u1_u12_u2_n171 ) );
  INV_X1 u1_u12_u2_U16 (.A( u1_u12_u2_n156 ) , .ZN( u1_u12_u2_n171 ) );
  INV_X1 u1_u12_u2_U17 (.A( u1_u12_u2_n120 ) , .ZN( u1_u12_u2_n188 ) );
  NAND2_X1 u1_u12_u2_U18 (.A2( u1_u12_u2_n122 ) , .ZN( u1_u12_u2_n150 ) , .A1( u1_u12_u2_n152 ) );
  INV_X1 u1_u12_u2_U19 (.A( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n170 ) );
  INV_X1 u1_u12_u2_U20 (.A( u1_u12_u2_n137 ) , .ZN( u1_u12_u2_n173 ) );
  NAND2_X1 u1_u12_u2_U21 (.A1( u1_u12_u2_n132 ) , .A2( u1_u12_u2_n139 ) , .ZN( u1_u12_u2_n157 ) );
  INV_X1 u1_u12_u2_U22 (.A( u1_u12_u2_n113 ) , .ZN( u1_u12_u2_n178 ) );
  INV_X1 u1_u12_u2_U23 (.A( u1_u12_u2_n139 ) , .ZN( u1_u12_u2_n175 ) );
  INV_X1 u1_u12_u2_U24 (.A( u1_u12_u2_n155 ) , .ZN( u1_u12_u2_n181 ) );
  INV_X1 u1_u12_u2_U25 (.A( u1_u12_u2_n119 ) , .ZN( u1_u12_u2_n177 ) );
  INV_X1 u1_u12_u2_U26 (.A( u1_u12_u2_n116 ) , .ZN( u1_u12_u2_n180 ) );
  INV_X1 u1_u12_u2_U27 (.A( u1_u12_u2_n131 ) , .ZN( u1_u12_u2_n179 ) );
  INV_X1 u1_u12_u2_U28 (.A( u1_u12_u2_n154 ) , .ZN( u1_u12_u2_n176 ) );
  NAND2_X1 u1_u12_u2_U29 (.A2( u1_u12_u2_n116 ) , .A1( u1_u12_u2_n117 ) , .ZN( u1_u12_u2_n118 ) );
  NOR2_X1 u1_u12_u2_U3 (.ZN( u1_u12_u2_n121 ) , .A2( u1_u12_u2_n177 ) , .A1( u1_u12_u2_n180 ) );
  INV_X1 u1_u12_u2_U30 (.A( u1_u12_u2_n132 ) , .ZN( u1_u12_u2_n182 ) );
  INV_X1 u1_u12_u2_U31 (.A( u1_u12_u2_n158 ) , .ZN( u1_u12_u2_n183 ) );
  OAI21_X1 u1_u12_u2_U32 (.A( u1_u12_u2_n156 ) , .B1( u1_u12_u2_n157 ) , .ZN( u1_u12_u2_n158 ) , .B2( u1_u12_u2_n179 ) );
  NOR2_X1 u1_u12_u2_U33 (.ZN( u1_u12_u2_n156 ) , .A1( u1_u12_u2_n166 ) , .A2( u1_u12_u2_n169 ) );
  NOR2_X1 u1_u12_u2_U34 (.A2( u1_u12_u2_n114 ) , .ZN( u1_u12_u2_n137 ) , .A1( u1_u12_u2_n140 ) );
  NOR2_X1 u1_u12_u2_U35 (.A2( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n153 ) , .A1( u1_u12_u2_n156 ) );
  AOI211_X1 u1_u12_u2_U36 (.ZN( u1_u12_u2_n130 ) , .C1( u1_u12_u2_n138 ) , .C2( u1_u12_u2_n179 ) , .B( u1_u12_u2_n96 ) , .A( u1_u12_u2_n97 ) );
  OAI22_X1 u1_u12_u2_U37 (.B1( u1_u12_u2_n133 ) , .A2( u1_u12_u2_n137 ) , .A1( u1_u12_u2_n152 ) , .B2( u1_u12_u2_n168 ) , .ZN( u1_u12_u2_n97 ) );
  OAI221_X1 u1_u12_u2_U38 (.B1( u1_u12_u2_n113 ) , .C1( u1_u12_u2_n132 ) , .A( u1_u12_u2_n149 ) , .B2( u1_u12_u2_n171 ) , .C2( u1_u12_u2_n172 ) , .ZN( u1_u12_u2_n96 ) );
  OAI221_X1 u1_u12_u2_U39 (.A( u1_u12_u2_n115 ) , .C2( u1_u12_u2_n123 ) , .B2( u1_u12_u2_n143 ) , .B1( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n163 ) , .C1( u1_u12_u2_n168 ) );
  INV_X1 u1_u12_u2_U4 (.A( u1_u12_u2_n134 ) , .ZN( u1_u12_u2_n185 ) );
  OAI21_X1 u1_u12_u2_U40 (.A( u1_u12_u2_n114 ) , .ZN( u1_u12_u2_n115 ) , .B1( u1_u12_u2_n176 ) , .B2( u1_u12_u2_n178 ) );
  OAI221_X1 u1_u12_u2_U41 (.A( u1_u12_u2_n135 ) , .B2( u1_u12_u2_n136 ) , .B1( u1_u12_u2_n137 ) , .ZN( u1_u12_u2_n162 ) , .C2( u1_u12_u2_n167 ) , .C1( u1_u12_u2_n185 ) );
  AND3_X1 u1_u12_u2_U42 (.A3( u1_u12_u2_n131 ) , .A2( u1_u12_u2_n132 ) , .A1( u1_u12_u2_n133 ) , .ZN( u1_u12_u2_n136 ) );
  AOI22_X1 u1_u12_u2_U43 (.ZN( u1_u12_u2_n135 ) , .B1( u1_u12_u2_n140 ) , .A1( u1_u12_u2_n156 ) , .B2( u1_u12_u2_n180 ) , .A2( u1_u12_u2_n188 ) );
  AOI21_X1 u1_u12_u2_U44 (.ZN( u1_u12_u2_n149 ) , .B1( u1_u12_u2_n173 ) , .B2( u1_u12_u2_n188 ) , .A( u1_u12_u2_n95 ) );
  AND3_X1 u1_u12_u2_U45 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n104 ) , .A3( u1_u12_u2_n156 ) , .ZN( u1_u12_u2_n95 ) );
  OAI21_X1 u1_u12_u2_U46 (.A( u1_u12_u2_n101 ) , .B2( u1_u12_u2_n121 ) , .B1( u1_u12_u2_n153 ) , .ZN( u1_u12_u2_n164 ) );
  NAND2_X1 u1_u12_u2_U47 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n107 ) , .ZN( u1_u12_u2_n155 ) );
  NAND2_X1 u1_u12_u2_U48 (.A2( u1_u12_u2_n105 ) , .A1( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n143 ) );
  NAND2_X1 u1_u12_u2_U49 (.A1( u1_u12_u2_n104 ) , .A2( u1_u12_u2_n106 ) , .ZN( u1_u12_u2_n152 ) );
  NOR4_X1 u1_u12_u2_U5 (.A4( u1_u12_u2_n124 ) , .A3( u1_u12_u2_n125 ) , .A2( u1_u12_u2_n126 ) , .A1( u1_u12_u2_n127 ) , .ZN( u1_u12_u2_n128 ) );
  NAND2_X1 u1_u12_u2_U50 (.A1( u1_u12_u2_n100 ) , .A2( u1_u12_u2_n105 ) , .ZN( u1_u12_u2_n132 ) );
  INV_X1 u1_u12_u2_U51 (.A( u1_u12_u2_n140 ) , .ZN( u1_u12_u2_n168 ) );
  INV_X1 u1_u12_u2_U52 (.A( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n167 ) );
  OAI21_X1 u1_u12_u2_U53 (.A( u1_u12_u2_n141 ) , .B2( u1_u12_u2_n142 ) , .ZN( u1_u12_u2_n146 ) , .B1( u1_u12_u2_n153 ) );
  OAI21_X1 u1_u12_u2_U54 (.A( u1_u12_u2_n140 ) , .ZN( u1_u12_u2_n141 ) , .B1( u1_u12_u2_n176 ) , .B2( u1_u12_u2_n177 ) );
  NOR3_X1 u1_u12_u2_U55 (.ZN( u1_u12_u2_n142 ) , .A3( u1_u12_u2_n175 ) , .A2( u1_u12_u2_n178 ) , .A1( u1_u12_u2_n181 ) );
  NAND2_X1 u1_u12_u2_U56 (.A1( u1_u12_u2_n102 ) , .A2( u1_u12_u2_n106 ) , .ZN( u1_u12_u2_n113 ) );
  NAND2_X1 u1_u12_u2_U57 (.A1( u1_u12_u2_n106 ) , .A2( u1_u12_u2_n107 ) , .ZN( u1_u12_u2_n131 ) );
  NAND2_X1 u1_u12_u2_U58 (.A1( u1_u12_u2_n103 ) , .A2( u1_u12_u2_n107 ) , .ZN( u1_u12_u2_n139 ) );
  NAND2_X1 u1_u12_u2_U59 (.A1( u1_u12_u2_n103 ) , .A2( u1_u12_u2_n105 ) , .ZN( u1_u12_u2_n133 ) );
  AOI21_X1 u1_u12_u2_U6 (.B2( u1_u12_u2_n119 ) , .ZN( u1_u12_u2_n127 ) , .A( u1_u12_u2_n137 ) , .B1( u1_u12_u2_n155 ) );
  NAND2_X1 u1_u12_u2_U60 (.A1( u1_u12_u2_n102 ) , .A2( u1_u12_u2_n103 ) , .ZN( u1_u12_u2_n154 ) );
  NAND2_X1 u1_u12_u2_U61 (.A2( u1_u12_u2_n103 ) , .A1( u1_u12_u2_n104 ) , .ZN( u1_u12_u2_n119 ) );
  NAND2_X1 u1_u12_u2_U62 (.A2( u1_u12_u2_n107 ) , .A1( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n123 ) );
  NAND2_X1 u1_u12_u2_U63 (.A1( u1_u12_u2_n104 ) , .A2( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n122 ) );
  INV_X1 u1_u12_u2_U64 (.A( u1_u12_u2_n114 ) , .ZN( u1_u12_u2_n172 ) );
  NAND2_X1 u1_u12_u2_U65 (.A2( u1_u12_u2_n100 ) , .A1( u1_u12_u2_n102 ) , .ZN( u1_u12_u2_n116 ) );
  NAND2_X1 u1_u12_u2_U66 (.A1( u1_u12_u2_n102 ) , .A2( u1_u12_u2_n108 ) , .ZN( u1_u12_u2_n120 ) );
  NAND2_X1 u1_u12_u2_U67 (.A2( u1_u12_u2_n105 ) , .A1( u1_u12_u2_n106 ) , .ZN( u1_u12_u2_n117 ) );
  INV_X1 u1_u12_u2_U68 (.ZN( u1_u12_u2_n187 ) , .A( u1_u12_u2_n99 ) );
  OAI21_X1 u1_u12_u2_U69 (.B1( u1_u12_u2_n137 ) , .B2( u1_u12_u2_n143 ) , .A( u1_u12_u2_n98 ) , .ZN( u1_u12_u2_n99 ) );
  AOI21_X1 u1_u12_u2_U7 (.ZN( u1_u12_u2_n124 ) , .B1( u1_u12_u2_n131 ) , .B2( u1_u12_u2_n143 ) , .A( u1_u12_u2_n172 ) );
  NOR2_X1 u1_u12_u2_U70 (.A2( u1_u12_X_16 ) , .ZN( u1_u12_u2_n140 ) , .A1( u1_u12_u2_n166 ) );
  NOR2_X1 u1_u12_u2_U71 (.A2( u1_u12_X_13 ) , .A1( u1_u12_X_14 ) , .ZN( u1_u12_u2_n100 ) );
  NOR2_X1 u1_u12_u2_U72 (.A2( u1_u12_X_16 ) , .A1( u1_u12_X_17 ) , .ZN( u1_u12_u2_n138 ) );
  NOR2_X1 u1_u12_u2_U73 (.A2( u1_u12_X_15 ) , .A1( u1_u12_X_18 ) , .ZN( u1_u12_u2_n104 ) );
  NOR2_X1 u1_u12_u2_U74 (.A2( u1_u12_X_14 ) , .ZN( u1_u12_u2_n103 ) , .A1( u1_u12_u2_n174 ) );
  NOR2_X1 u1_u12_u2_U75 (.A2( u1_u12_X_15 ) , .ZN( u1_u12_u2_n102 ) , .A1( u1_u12_u2_n165 ) );
  NOR2_X1 u1_u12_u2_U76 (.A2( u1_u12_X_17 ) , .ZN( u1_u12_u2_n114 ) , .A1( u1_u12_u2_n169 ) );
  AND2_X1 u1_u12_u2_U77 (.A1( u1_u12_X_15 ) , .ZN( u1_u12_u2_n105 ) , .A2( u1_u12_u2_n165 ) );
  AND2_X1 u1_u12_u2_U78 (.A2( u1_u12_X_15 ) , .A1( u1_u12_X_18 ) , .ZN( u1_u12_u2_n107 ) );
  AND2_X1 u1_u12_u2_U79 (.A1( u1_u12_X_14 ) , .ZN( u1_u12_u2_n106 ) , .A2( u1_u12_u2_n174 ) );
  AOI21_X1 u1_u12_u2_U8 (.B2( u1_u12_u2_n120 ) , .B1( u1_u12_u2_n121 ) , .ZN( u1_u12_u2_n126 ) , .A( u1_u12_u2_n167 ) );
  AND2_X1 u1_u12_u2_U80 (.A1( u1_u12_X_13 ) , .A2( u1_u12_X_14 ) , .ZN( u1_u12_u2_n108 ) );
  INV_X1 u1_u12_u2_U81 (.A( u1_u12_X_16 ) , .ZN( u1_u12_u2_n169 ) );
  INV_X1 u1_u12_u2_U82 (.A( u1_u12_X_17 ) , .ZN( u1_u12_u2_n166 ) );
  INV_X1 u1_u12_u2_U83 (.A( u1_u12_X_13 ) , .ZN( u1_u12_u2_n174 ) );
  INV_X1 u1_u12_u2_U84 (.A( u1_u12_X_18 ) , .ZN( u1_u12_u2_n165 ) );
  NAND4_X1 u1_u12_u2_U85 (.ZN( u1_out12_30 ) , .A4( u1_u12_u2_n147 ) , .A3( u1_u12_u2_n148 ) , .A2( u1_u12_u2_n149 ) , .A1( u1_u12_u2_n187 ) );
  AOI21_X1 u1_u12_u2_U86 (.B2( u1_u12_u2_n138 ) , .ZN( u1_u12_u2_n148 ) , .A( u1_u12_u2_n162 ) , .B1( u1_u12_u2_n182 ) );
  NOR3_X1 u1_u12_u2_U87 (.A3( u1_u12_u2_n144 ) , .A2( u1_u12_u2_n145 ) , .A1( u1_u12_u2_n146 ) , .ZN( u1_u12_u2_n147 ) );
  NAND4_X1 u1_u12_u2_U88 (.ZN( u1_out12_24 ) , .A4( u1_u12_u2_n111 ) , .A3( u1_u12_u2_n112 ) , .A1( u1_u12_u2_n130 ) , .A2( u1_u12_u2_n187 ) );
  AOI221_X1 u1_u12_u2_U89 (.A( u1_u12_u2_n109 ) , .B1( u1_u12_u2_n110 ) , .ZN( u1_u12_u2_n111 ) , .C1( u1_u12_u2_n134 ) , .C2( u1_u12_u2_n170 ) , .B2( u1_u12_u2_n173 ) );
  OAI22_X1 u1_u12_u2_U9 (.ZN( u1_u12_u2_n109 ) , .A2( u1_u12_u2_n113 ) , .B2( u1_u12_u2_n133 ) , .B1( u1_u12_u2_n167 ) , .A1( u1_u12_u2_n168 ) );
  AOI21_X1 u1_u12_u2_U90 (.ZN( u1_u12_u2_n112 ) , .B2( u1_u12_u2_n156 ) , .A( u1_u12_u2_n164 ) , .B1( u1_u12_u2_n181 ) );
  NAND4_X1 u1_u12_u2_U91 (.ZN( u1_out12_16 ) , .A4( u1_u12_u2_n128 ) , .A3( u1_u12_u2_n129 ) , .A1( u1_u12_u2_n130 ) , .A2( u1_u12_u2_n186 ) );
  AOI22_X1 u1_u12_u2_U92 (.A2( u1_u12_u2_n118 ) , .ZN( u1_u12_u2_n129 ) , .A1( u1_u12_u2_n140 ) , .B1( u1_u12_u2_n157 ) , .B2( u1_u12_u2_n170 ) );
  INV_X1 u1_u12_u2_U93 (.A( u1_u12_u2_n163 ) , .ZN( u1_u12_u2_n186 ) );
  OR4_X1 u1_u12_u2_U94 (.ZN( u1_out12_6 ) , .A4( u1_u12_u2_n161 ) , .A3( u1_u12_u2_n162 ) , .A2( u1_u12_u2_n163 ) , .A1( u1_u12_u2_n164 ) );
  OR3_X1 u1_u12_u2_U95 (.A2( u1_u12_u2_n159 ) , .A1( u1_u12_u2_n160 ) , .ZN( u1_u12_u2_n161 ) , .A3( u1_u12_u2_n183 ) );
  AOI21_X1 u1_u12_u2_U96 (.B2( u1_u12_u2_n154 ) , .B1( u1_u12_u2_n155 ) , .ZN( u1_u12_u2_n159 ) , .A( u1_u12_u2_n167 ) );
  NAND3_X1 u1_u12_u2_U97 (.A2( u1_u12_u2_n117 ) , .A1( u1_u12_u2_n122 ) , .A3( u1_u12_u2_n123 ) , .ZN( u1_u12_u2_n134 ) );
  NAND3_X1 u1_u12_u2_U98 (.ZN( u1_u12_u2_n110 ) , .A2( u1_u12_u2_n131 ) , .A3( u1_u12_u2_n139 ) , .A1( u1_u12_u2_n154 ) );
  NAND3_X1 u1_u12_u2_U99 (.A2( u1_u12_u2_n100 ) , .ZN( u1_u12_u2_n101 ) , .A1( u1_u12_u2_n104 ) , .A3( u1_u12_u2_n114 ) );
  AOI22_X1 u1_u12_u6_U10 (.A2( u1_u12_u6_n151 ) , .B2( u1_u12_u6_n161 ) , .A1( u1_u12_u6_n167 ) , .B1( u1_u12_u6_n170 ) , .ZN( u1_u12_u6_n89 ) );
  AOI21_X1 u1_u12_u6_U11 (.B1( u1_u12_u6_n107 ) , .B2( u1_u12_u6_n132 ) , .A( u1_u12_u6_n158 ) , .ZN( u1_u12_u6_n88 ) );
  AOI21_X1 u1_u12_u6_U12 (.B2( u1_u12_u6_n147 ) , .B1( u1_u12_u6_n148 ) , .ZN( u1_u12_u6_n149 ) , .A( u1_u12_u6_n158 ) );
  AOI21_X1 u1_u12_u6_U13 (.ZN( u1_u12_u6_n106 ) , .A( u1_u12_u6_n142 ) , .B2( u1_u12_u6_n159 ) , .B1( u1_u12_u6_n164 ) );
  INV_X1 u1_u12_u6_U14 (.A( u1_u12_u6_n155 ) , .ZN( u1_u12_u6_n161 ) );
  INV_X1 u1_u12_u6_U15 (.A( u1_u12_u6_n128 ) , .ZN( u1_u12_u6_n164 ) );
  NAND2_X1 u1_u12_u6_U16 (.ZN( u1_u12_u6_n110 ) , .A1( u1_u12_u6_n122 ) , .A2( u1_u12_u6_n129 ) );
  NAND2_X1 u1_u12_u6_U17 (.ZN( u1_u12_u6_n124 ) , .A2( u1_u12_u6_n146 ) , .A1( u1_u12_u6_n148 ) );
  INV_X1 u1_u12_u6_U18 (.A( u1_u12_u6_n132 ) , .ZN( u1_u12_u6_n171 ) );
  AND2_X1 u1_u12_u6_U19 (.A1( u1_u12_u6_n100 ) , .ZN( u1_u12_u6_n130 ) , .A2( u1_u12_u6_n147 ) );
  INV_X1 u1_u12_u6_U20 (.A( u1_u12_u6_n127 ) , .ZN( u1_u12_u6_n173 ) );
  INV_X1 u1_u12_u6_U21 (.A( u1_u12_u6_n121 ) , .ZN( u1_u12_u6_n167 ) );
  INV_X1 u1_u12_u6_U22 (.A( u1_u12_u6_n100 ) , .ZN( u1_u12_u6_n169 ) );
  INV_X1 u1_u12_u6_U23 (.A( u1_u12_u6_n123 ) , .ZN( u1_u12_u6_n170 ) );
  INV_X1 u1_u12_u6_U24 (.A( u1_u12_u6_n113 ) , .ZN( u1_u12_u6_n168 ) );
  AND2_X1 u1_u12_u6_U25 (.A1( u1_u12_u6_n107 ) , .A2( u1_u12_u6_n119 ) , .ZN( u1_u12_u6_n133 ) );
  AND2_X1 u1_u12_u6_U26 (.A2( u1_u12_u6_n121 ) , .A1( u1_u12_u6_n122 ) , .ZN( u1_u12_u6_n131 ) );
  AND3_X1 u1_u12_u6_U27 (.ZN( u1_u12_u6_n120 ) , .A2( u1_u12_u6_n127 ) , .A1( u1_u12_u6_n132 ) , .A3( u1_u12_u6_n145 ) );
  INV_X1 u1_u12_u6_U28 (.A( u1_u12_u6_n146 ) , .ZN( u1_u12_u6_n163 ) );
  AOI222_X1 u1_u12_u6_U29 (.ZN( u1_u12_u6_n114 ) , .A1( u1_u12_u6_n118 ) , .A2( u1_u12_u6_n126 ) , .B2( u1_u12_u6_n151 ) , .C2( u1_u12_u6_n159 ) , .C1( u1_u12_u6_n168 ) , .B1( u1_u12_u6_n169 ) );
  INV_X1 u1_u12_u6_U3 (.A( u1_u12_u6_n110 ) , .ZN( u1_u12_u6_n166 ) );
  NOR2_X1 u1_u12_u6_U30 (.A1( u1_u12_u6_n162 ) , .A2( u1_u12_u6_n165 ) , .ZN( u1_u12_u6_n98 ) );
  AOI211_X1 u1_u12_u6_U31 (.B( u1_u12_u6_n134 ) , .A( u1_u12_u6_n135 ) , .C1( u1_u12_u6_n136 ) , .ZN( u1_u12_u6_n137 ) , .C2( u1_u12_u6_n151 ) );
  AOI21_X1 u1_u12_u6_U32 (.B2( u1_u12_u6_n132 ) , .B1( u1_u12_u6_n133 ) , .ZN( u1_u12_u6_n134 ) , .A( u1_u12_u6_n158 ) );
  AOI21_X1 u1_u12_u6_U33 (.B1( u1_u12_u6_n131 ) , .ZN( u1_u12_u6_n135 ) , .A( u1_u12_u6_n144 ) , .B2( u1_u12_u6_n146 ) );
  NAND4_X1 u1_u12_u6_U34 (.A4( u1_u12_u6_n127 ) , .A3( u1_u12_u6_n128 ) , .A2( u1_u12_u6_n129 ) , .A1( u1_u12_u6_n130 ) , .ZN( u1_u12_u6_n136 ) );
  NAND2_X1 u1_u12_u6_U35 (.A1( u1_u12_u6_n144 ) , .ZN( u1_u12_u6_n151 ) , .A2( u1_u12_u6_n158 ) );
  NAND2_X1 u1_u12_u6_U36 (.ZN( u1_u12_u6_n132 ) , .A1( u1_u12_u6_n91 ) , .A2( u1_u12_u6_n97 ) );
  AOI22_X1 u1_u12_u6_U37 (.B2( u1_u12_u6_n110 ) , .B1( u1_u12_u6_n111 ) , .A1( u1_u12_u6_n112 ) , .ZN( u1_u12_u6_n115 ) , .A2( u1_u12_u6_n161 ) );
  NAND4_X1 u1_u12_u6_U38 (.A3( u1_u12_u6_n109 ) , .ZN( u1_u12_u6_n112 ) , .A4( u1_u12_u6_n132 ) , .A2( u1_u12_u6_n147 ) , .A1( u1_u12_u6_n166 ) );
  NOR2_X1 u1_u12_u6_U39 (.ZN( u1_u12_u6_n109 ) , .A1( u1_u12_u6_n170 ) , .A2( u1_u12_u6_n173 ) );
  INV_X1 u1_u12_u6_U4 (.A( u1_u12_u6_n142 ) , .ZN( u1_u12_u6_n174 ) );
  NOR2_X1 u1_u12_u6_U40 (.A2( u1_u12_u6_n126 ) , .ZN( u1_u12_u6_n155 ) , .A1( u1_u12_u6_n160 ) );
  NAND2_X1 u1_u12_u6_U41 (.ZN( u1_u12_u6_n146 ) , .A2( u1_u12_u6_n94 ) , .A1( u1_u12_u6_n99 ) );
  AOI21_X1 u1_u12_u6_U42 (.A( u1_u12_u6_n144 ) , .B2( u1_u12_u6_n145 ) , .B1( u1_u12_u6_n146 ) , .ZN( u1_u12_u6_n150 ) );
  INV_X1 u1_u12_u6_U43 (.A( u1_u12_u6_n111 ) , .ZN( u1_u12_u6_n158 ) );
  NAND2_X1 u1_u12_u6_U44 (.ZN( u1_u12_u6_n127 ) , .A1( u1_u12_u6_n91 ) , .A2( u1_u12_u6_n92 ) );
  NAND2_X1 u1_u12_u6_U45 (.ZN( u1_u12_u6_n129 ) , .A2( u1_u12_u6_n95 ) , .A1( u1_u12_u6_n96 ) );
  INV_X1 u1_u12_u6_U46 (.A( u1_u12_u6_n144 ) , .ZN( u1_u12_u6_n159 ) );
  NAND2_X1 u1_u12_u6_U47 (.ZN( u1_u12_u6_n145 ) , .A2( u1_u12_u6_n97 ) , .A1( u1_u12_u6_n98 ) );
  NAND2_X1 u1_u12_u6_U48 (.ZN( u1_u12_u6_n148 ) , .A2( u1_u12_u6_n92 ) , .A1( u1_u12_u6_n94 ) );
  NAND2_X1 u1_u12_u6_U49 (.ZN( u1_u12_u6_n108 ) , .A2( u1_u12_u6_n139 ) , .A1( u1_u12_u6_n144 ) );
  NAND2_X1 u1_u12_u6_U5 (.A2( u1_u12_u6_n143 ) , .ZN( u1_u12_u6_n152 ) , .A1( u1_u12_u6_n166 ) );
  NAND2_X1 u1_u12_u6_U50 (.ZN( u1_u12_u6_n121 ) , .A2( u1_u12_u6_n95 ) , .A1( u1_u12_u6_n97 ) );
  NAND2_X1 u1_u12_u6_U51 (.ZN( u1_u12_u6_n107 ) , .A2( u1_u12_u6_n92 ) , .A1( u1_u12_u6_n95 ) );
  AND2_X1 u1_u12_u6_U52 (.ZN( u1_u12_u6_n118 ) , .A2( u1_u12_u6_n91 ) , .A1( u1_u12_u6_n99 ) );
  NAND2_X1 u1_u12_u6_U53 (.ZN( u1_u12_u6_n147 ) , .A2( u1_u12_u6_n98 ) , .A1( u1_u12_u6_n99 ) );
  NAND2_X1 u1_u12_u6_U54 (.ZN( u1_u12_u6_n128 ) , .A1( u1_u12_u6_n94 ) , .A2( u1_u12_u6_n96 ) );
  NAND2_X1 u1_u12_u6_U55 (.ZN( u1_u12_u6_n119 ) , .A2( u1_u12_u6_n95 ) , .A1( u1_u12_u6_n99 ) );
  NAND2_X1 u1_u12_u6_U56 (.ZN( u1_u12_u6_n123 ) , .A2( u1_u12_u6_n91 ) , .A1( u1_u12_u6_n96 ) );
  NAND2_X1 u1_u12_u6_U57 (.ZN( u1_u12_u6_n100 ) , .A2( u1_u12_u6_n92 ) , .A1( u1_u12_u6_n98 ) );
  NAND2_X1 u1_u12_u6_U58 (.ZN( u1_u12_u6_n122 ) , .A1( u1_u12_u6_n94 ) , .A2( u1_u12_u6_n97 ) );
  INV_X1 u1_u12_u6_U59 (.A( u1_u12_u6_n139 ) , .ZN( u1_u12_u6_n160 ) );
  AOI22_X1 u1_u12_u6_U6 (.B2( u1_u12_u6_n101 ) , .A1( u1_u12_u6_n102 ) , .ZN( u1_u12_u6_n103 ) , .B1( u1_u12_u6_n160 ) , .A2( u1_u12_u6_n161 ) );
  NAND2_X1 u1_u12_u6_U60 (.ZN( u1_u12_u6_n113 ) , .A1( u1_u12_u6_n96 ) , .A2( u1_u12_u6_n98 ) );
  NOR2_X1 u1_u12_u6_U61 (.A2( u1_u12_X_40 ) , .A1( u1_u12_X_41 ) , .ZN( u1_u12_u6_n126 ) );
  NOR2_X1 u1_u12_u6_U62 (.A2( u1_u12_X_39 ) , .A1( u1_u12_X_42 ) , .ZN( u1_u12_u6_n92 ) );
  NOR2_X1 u1_u12_u6_U63 (.A2( u1_u12_X_39 ) , .A1( u1_u12_u6_n156 ) , .ZN( u1_u12_u6_n97 ) );
  NOR2_X1 u1_u12_u6_U64 (.A2( u1_u12_X_38 ) , .A1( u1_u12_u6_n165 ) , .ZN( u1_u12_u6_n95 ) );
  NOR2_X1 u1_u12_u6_U65 (.A2( u1_u12_X_41 ) , .ZN( u1_u12_u6_n111 ) , .A1( u1_u12_u6_n157 ) );
  NOR2_X1 u1_u12_u6_U66 (.A2( u1_u12_X_37 ) , .A1( u1_u12_u6_n162 ) , .ZN( u1_u12_u6_n94 ) );
  NOR2_X1 u1_u12_u6_U67 (.A2( u1_u12_X_37 ) , .A1( u1_u12_X_38 ) , .ZN( u1_u12_u6_n91 ) );
  NAND2_X1 u1_u12_u6_U68 (.A1( u1_u12_X_41 ) , .ZN( u1_u12_u6_n144 ) , .A2( u1_u12_u6_n157 ) );
  NAND2_X1 u1_u12_u6_U69 (.A2( u1_u12_X_40 ) , .A1( u1_u12_X_41 ) , .ZN( u1_u12_u6_n139 ) );
  NOR2_X1 u1_u12_u6_U7 (.A1( u1_u12_u6_n118 ) , .ZN( u1_u12_u6_n143 ) , .A2( u1_u12_u6_n168 ) );
  AND2_X1 u1_u12_u6_U70 (.A1( u1_u12_X_39 ) , .A2( u1_u12_u6_n156 ) , .ZN( u1_u12_u6_n96 ) );
  AND2_X1 u1_u12_u6_U71 (.A1( u1_u12_X_39 ) , .A2( u1_u12_X_42 ) , .ZN( u1_u12_u6_n99 ) );
  INV_X1 u1_u12_u6_U72 (.A( u1_u12_X_40 ) , .ZN( u1_u12_u6_n157 ) );
  INV_X1 u1_u12_u6_U73 (.A( u1_u12_X_37 ) , .ZN( u1_u12_u6_n165 ) );
  INV_X1 u1_u12_u6_U74 (.A( u1_u12_X_38 ) , .ZN( u1_u12_u6_n162 ) );
  INV_X1 u1_u12_u6_U75 (.A( u1_u12_X_42 ) , .ZN( u1_u12_u6_n156 ) );
  NAND4_X1 u1_u12_u6_U76 (.ZN( u1_out12_32 ) , .A4( u1_u12_u6_n103 ) , .A3( u1_u12_u6_n104 ) , .A2( u1_u12_u6_n105 ) , .A1( u1_u12_u6_n106 ) );
  AOI22_X1 u1_u12_u6_U77 (.ZN( u1_u12_u6_n105 ) , .A2( u1_u12_u6_n108 ) , .A1( u1_u12_u6_n118 ) , .B2( u1_u12_u6_n126 ) , .B1( u1_u12_u6_n171 ) );
  AOI22_X1 u1_u12_u6_U78 (.ZN( u1_u12_u6_n104 ) , .A1( u1_u12_u6_n111 ) , .B1( u1_u12_u6_n124 ) , .B2( u1_u12_u6_n151 ) , .A2( u1_u12_u6_n93 ) );
  NAND4_X1 u1_u12_u6_U79 (.ZN( u1_out12_12 ) , .A4( u1_u12_u6_n114 ) , .A3( u1_u12_u6_n115 ) , .A2( u1_u12_u6_n116 ) , .A1( u1_u12_u6_n117 ) );
  INV_X1 u1_u12_u6_U8 (.ZN( u1_u12_u6_n172 ) , .A( u1_u12_u6_n88 ) );
  OAI22_X1 u1_u12_u6_U80 (.B2( u1_u12_u6_n111 ) , .ZN( u1_u12_u6_n116 ) , .B1( u1_u12_u6_n126 ) , .A2( u1_u12_u6_n164 ) , .A1( u1_u12_u6_n167 ) );
  OAI21_X1 u1_u12_u6_U81 (.A( u1_u12_u6_n108 ) , .ZN( u1_u12_u6_n117 ) , .B2( u1_u12_u6_n141 ) , .B1( u1_u12_u6_n163 ) );
  OAI211_X1 u1_u12_u6_U82 (.ZN( u1_out12_22 ) , .B( u1_u12_u6_n137 ) , .A( u1_u12_u6_n138 ) , .C2( u1_u12_u6_n139 ) , .C1( u1_u12_u6_n140 ) );
  AOI22_X1 u1_u12_u6_U83 (.B1( u1_u12_u6_n124 ) , .A2( u1_u12_u6_n125 ) , .A1( u1_u12_u6_n126 ) , .ZN( u1_u12_u6_n138 ) , .B2( u1_u12_u6_n161 ) );
  AND4_X1 u1_u12_u6_U84 (.A3( u1_u12_u6_n119 ) , .A1( u1_u12_u6_n120 ) , .A4( u1_u12_u6_n129 ) , .ZN( u1_u12_u6_n140 ) , .A2( u1_u12_u6_n143 ) );
  OAI211_X1 u1_u12_u6_U85 (.ZN( u1_out12_7 ) , .B( u1_u12_u6_n153 ) , .C2( u1_u12_u6_n154 ) , .C1( u1_u12_u6_n155 ) , .A( u1_u12_u6_n174 ) );
  NOR3_X1 u1_u12_u6_U86 (.A1( u1_u12_u6_n141 ) , .ZN( u1_u12_u6_n154 ) , .A3( u1_u12_u6_n164 ) , .A2( u1_u12_u6_n171 ) );
  AOI211_X1 u1_u12_u6_U87 (.B( u1_u12_u6_n149 ) , .A( u1_u12_u6_n150 ) , .C2( u1_u12_u6_n151 ) , .C1( u1_u12_u6_n152 ) , .ZN( u1_u12_u6_n153 ) );
  NAND3_X1 u1_u12_u6_U88 (.A2( u1_u12_u6_n123 ) , .ZN( u1_u12_u6_n125 ) , .A1( u1_u12_u6_n130 ) , .A3( u1_u12_u6_n131 ) );
  NAND3_X1 u1_u12_u6_U89 (.A3( u1_u12_u6_n133 ) , .ZN( u1_u12_u6_n141 ) , .A1( u1_u12_u6_n145 ) , .A2( u1_u12_u6_n148 ) );
  OAI21_X1 u1_u12_u6_U9 (.A( u1_u12_u6_n159 ) , .B1( u1_u12_u6_n169 ) , .B2( u1_u12_u6_n173 ) , .ZN( u1_u12_u6_n90 ) );
  NAND3_X1 u1_u12_u6_U90 (.ZN( u1_u12_u6_n101 ) , .A3( u1_u12_u6_n107 ) , .A2( u1_u12_u6_n121 ) , .A1( u1_u12_u6_n127 ) );
  NAND3_X1 u1_u12_u6_U91 (.ZN( u1_u12_u6_n102 ) , .A3( u1_u12_u6_n130 ) , .A2( u1_u12_u6_n145 ) , .A1( u1_u12_u6_n166 ) );
  NAND3_X1 u1_u12_u6_U92 (.A3( u1_u12_u6_n113 ) , .A1( u1_u12_u6_n119 ) , .A2( u1_u12_u6_n123 ) , .ZN( u1_u12_u6_n93 ) );
  NAND3_X1 u1_u12_u6_U93 (.ZN( u1_u12_u6_n142 ) , .A2( u1_u12_u6_n172 ) , .A3( u1_u12_u6_n89 ) , .A1( u1_u12_u6_n90 ) );
  AND3_X1 u1_u12_u7_U10 (.A3( u1_u12_u7_n110 ) , .A2( u1_u12_u7_n127 ) , .A1( u1_u12_u7_n132 ) , .ZN( u1_u12_u7_n92 ) );
  OAI21_X1 u1_u12_u7_U11 (.A( u1_u12_u7_n161 ) , .B1( u1_u12_u7_n168 ) , .B2( u1_u12_u7_n173 ) , .ZN( u1_u12_u7_n91 ) );
  AOI211_X1 u1_u12_u7_U12 (.A( u1_u12_u7_n117 ) , .ZN( u1_u12_u7_n118 ) , .C2( u1_u12_u7_n126 ) , .C1( u1_u12_u7_n177 ) , .B( u1_u12_u7_n180 ) );
  OAI22_X1 u1_u12_u7_U13 (.B1( u1_u12_u7_n115 ) , .ZN( u1_u12_u7_n117 ) , .A2( u1_u12_u7_n133 ) , .A1( u1_u12_u7_n137 ) , .B2( u1_u12_u7_n162 ) );
  INV_X1 u1_u12_u7_U14 (.A( u1_u12_u7_n116 ) , .ZN( u1_u12_u7_n180 ) );
  NOR3_X1 u1_u12_u7_U15 (.ZN( u1_u12_u7_n115 ) , .A3( u1_u12_u7_n145 ) , .A2( u1_u12_u7_n168 ) , .A1( u1_u12_u7_n169 ) );
  OAI211_X1 u1_u12_u7_U16 (.B( u1_u12_u7_n122 ) , .A( u1_u12_u7_n123 ) , .C2( u1_u12_u7_n124 ) , .ZN( u1_u12_u7_n154 ) , .C1( u1_u12_u7_n162 ) );
  AOI222_X1 u1_u12_u7_U17 (.ZN( u1_u12_u7_n122 ) , .C2( u1_u12_u7_n126 ) , .C1( u1_u12_u7_n145 ) , .B1( u1_u12_u7_n161 ) , .A2( u1_u12_u7_n165 ) , .B2( u1_u12_u7_n170 ) , .A1( u1_u12_u7_n176 ) );
  INV_X1 u1_u12_u7_U18 (.A( u1_u12_u7_n133 ) , .ZN( u1_u12_u7_n176 ) );
  NOR3_X1 u1_u12_u7_U19 (.A2( u1_u12_u7_n134 ) , .A1( u1_u12_u7_n135 ) , .ZN( u1_u12_u7_n136 ) , .A3( u1_u12_u7_n171 ) );
  NOR2_X1 u1_u12_u7_U20 (.A1( u1_u12_u7_n130 ) , .A2( u1_u12_u7_n134 ) , .ZN( u1_u12_u7_n153 ) );
  INV_X1 u1_u12_u7_U21 (.A( u1_u12_u7_n101 ) , .ZN( u1_u12_u7_n165 ) );
  NOR2_X1 u1_u12_u7_U22 (.ZN( u1_u12_u7_n111 ) , .A2( u1_u12_u7_n134 ) , .A1( u1_u12_u7_n169 ) );
  AOI21_X1 u1_u12_u7_U23 (.ZN( u1_u12_u7_n104 ) , .B2( u1_u12_u7_n112 ) , .B1( u1_u12_u7_n127 ) , .A( u1_u12_u7_n164 ) );
  AOI21_X1 u1_u12_u7_U24 (.ZN( u1_u12_u7_n106 ) , .B1( u1_u12_u7_n133 ) , .B2( u1_u12_u7_n146 ) , .A( u1_u12_u7_n162 ) );
  AOI21_X1 u1_u12_u7_U25 (.A( u1_u12_u7_n101 ) , .ZN( u1_u12_u7_n107 ) , .B2( u1_u12_u7_n128 ) , .B1( u1_u12_u7_n175 ) );
  INV_X1 u1_u12_u7_U26 (.A( u1_u12_u7_n138 ) , .ZN( u1_u12_u7_n171 ) );
  INV_X1 u1_u12_u7_U27 (.A( u1_u12_u7_n131 ) , .ZN( u1_u12_u7_n177 ) );
  INV_X1 u1_u12_u7_U28 (.A( u1_u12_u7_n110 ) , .ZN( u1_u12_u7_n174 ) );
  NAND2_X1 u1_u12_u7_U29 (.A1( u1_u12_u7_n129 ) , .A2( u1_u12_u7_n132 ) , .ZN( u1_u12_u7_n149 ) );
  OAI21_X1 u1_u12_u7_U3 (.ZN( u1_u12_u7_n159 ) , .A( u1_u12_u7_n165 ) , .B2( u1_u12_u7_n171 ) , .B1( u1_u12_u7_n174 ) );
  NAND2_X1 u1_u12_u7_U30 (.A1( u1_u12_u7_n113 ) , .A2( u1_u12_u7_n124 ) , .ZN( u1_u12_u7_n130 ) );
  INV_X1 u1_u12_u7_U31 (.A( u1_u12_u7_n112 ) , .ZN( u1_u12_u7_n173 ) );
  INV_X1 u1_u12_u7_U32 (.A( u1_u12_u7_n128 ) , .ZN( u1_u12_u7_n168 ) );
  INV_X1 u1_u12_u7_U33 (.A( u1_u12_u7_n148 ) , .ZN( u1_u12_u7_n169 ) );
  INV_X1 u1_u12_u7_U34 (.A( u1_u12_u7_n127 ) , .ZN( u1_u12_u7_n179 ) );
  NOR2_X1 u1_u12_u7_U35 (.ZN( u1_u12_u7_n101 ) , .A2( u1_u12_u7_n150 ) , .A1( u1_u12_u7_n156 ) );
  AOI211_X1 u1_u12_u7_U36 (.B( u1_u12_u7_n154 ) , .A( u1_u12_u7_n155 ) , .C1( u1_u12_u7_n156 ) , .ZN( u1_u12_u7_n157 ) , .C2( u1_u12_u7_n172 ) );
  INV_X1 u1_u12_u7_U37 (.A( u1_u12_u7_n153 ) , .ZN( u1_u12_u7_n172 ) );
  AOI211_X1 u1_u12_u7_U38 (.B( u1_u12_u7_n139 ) , .A( u1_u12_u7_n140 ) , .C2( u1_u12_u7_n141 ) , .ZN( u1_u12_u7_n142 ) , .C1( u1_u12_u7_n156 ) );
  NAND4_X1 u1_u12_u7_U39 (.A3( u1_u12_u7_n127 ) , .A2( u1_u12_u7_n128 ) , .A1( u1_u12_u7_n129 ) , .ZN( u1_u12_u7_n141 ) , .A4( u1_u12_u7_n147 ) );
  INV_X1 u1_u12_u7_U4 (.A( u1_u12_u7_n111 ) , .ZN( u1_u12_u7_n170 ) );
  AOI21_X1 u1_u12_u7_U40 (.A( u1_u12_u7_n137 ) , .B1( u1_u12_u7_n138 ) , .ZN( u1_u12_u7_n139 ) , .B2( u1_u12_u7_n146 ) );
  OAI22_X1 u1_u12_u7_U41 (.B1( u1_u12_u7_n136 ) , .ZN( u1_u12_u7_n140 ) , .A1( u1_u12_u7_n153 ) , .B2( u1_u12_u7_n162 ) , .A2( u1_u12_u7_n164 ) );
  AOI21_X1 u1_u12_u7_U42 (.ZN( u1_u12_u7_n123 ) , .B1( u1_u12_u7_n165 ) , .B2( u1_u12_u7_n177 ) , .A( u1_u12_u7_n97 ) );
  AOI21_X1 u1_u12_u7_U43 (.B2( u1_u12_u7_n113 ) , .B1( u1_u12_u7_n124 ) , .A( u1_u12_u7_n125 ) , .ZN( u1_u12_u7_n97 ) );
  INV_X1 u1_u12_u7_U44 (.A( u1_u12_u7_n125 ) , .ZN( u1_u12_u7_n161 ) );
  INV_X1 u1_u12_u7_U45 (.A( u1_u12_u7_n152 ) , .ZN( u1_u12_u7_n162 ) );
  AOI22_X1 u1_u12_u7_U46 (.A2( u1_u12_u7_n114 ) , .ZN( u1_u12_u7_n119 ) , .B1( u1_u12_u7_n130 ) , .A1( u1_u12_u7_n156 ) , .B2( u1_u12_u7_n165 ) );
  NAND2_X1 u1_u12_u7_U47 (.A2( u1_u12_u7_n112 ) , .ZN( u1_u12_u7_n114 ) , .A1( u1_u12_u7_n175 ) );
  AND2_X1 u1_u12_u7_U48 (.ZN( u1_u12_u7_n145 ) , .A2( u1_u12_u7_n98 ) , .A1( u1_u12_u7_n99 ) );
  NOR2_X1 u1_u12_u7_U49 (.ZN( u1_u12_u7_n137 ) , .A1( u1_u12_u7_n150 ) , .A2( u1_u12_u7_n161 ) );
  INV_X1 u1_u12_u7_U5 (.A( u1_u12_u7_n149 ) , .ZN( u1_u12_u7_n175 ) );
  AOI21_X1 u1_u12_u7_U50 (.ZN( u1_u12_u7_n105 ) , .B2( u1_u12_u7_n110 ) , .A( u1_u12_u7_n125 ) , .B1( u1_u12_u7_n147 ) );
  NAND2_X1 u1_u12_u7_U51 (.ZN( u1_u12_u7_n146 ) , .A1( u1_u12_u7_n95 ) , .A2( u1_u12_u7_n98 ) );
  NAND2_X1 u1_u12_u7_U52 (.A2( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n147 ) , .A1( u1_u12_u7_n93 ) );
  NAND2_X1 u1_u12_u7_U53 (.A1( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n127 ) , .A2( u1_u12_u7_n99 ) );
  OR2_X1 u1_u12_u7_U54 (.ZN( u1_u12_u7_n126 ) , .A2( u1_u12_u7_n152 ) , .A1( u1_u12_u7_n156 ) );
  NAND2_X1 u1_u12_u7_U55 (.A2( u1_u12_u7_n102 ) , .A1( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n133 ) );
  NAND2_X1 u1_u12_u7_U56 (.ZN( u1_u12_u7_n112 ) , .A2( u1_u12_u7_n96 ) , .A1( u1_u12_u7_n99 ) );
  NAND2_X1 u1_u12_u7_U57 (.A2( u1_u12_u7_n102 ) , .ZN( u1_u12_u7_n128 ) , .A1( u1_u12_u7_n98 ) );
  NAND2_X1 u1_u12_u7_U58 (.A1( u1_u12_u7_n100 ) , .ZN( u1_u12_u7_n113 ) , .A2( u1_u12_u7_n93 ) );
  NAND2_X1 u1_u12_u7_U59 (.A2( u1_u12_u7_n102 ) , .ZN( u1_u12_u7_n124 ) , .A1( u1_u12_u7_n96 ) );
  INV_X1 u1_u12_u7_U6 (.A( u1_u12_u7_n154 ) , .ZN( u1_u12_u7_n178 ) );
  NAND2_X1 u1_u12_u7_U60 (.ZN( u1_u12_u7_n110 ) , .A1( u1_u12_u7_n95 ) , .A2( u1_u12_u7_n96 ) );
  INV_X1 u1_u12_u7_U61 (.A( u1_u12_u7_n150 ) , .ZN( u1_u12_u7_n164 ) );
  AND2_X1 u1_u12_u7_U62 (.ZN( u1_u12_u7_n134 ) , .A1( u1_u12_u7_n93 ) , .A2( u1_u12_u7_n98 ) );
  NAND2_X1 u1_u12_u7_U63 (.A1( u1_u12_u7_n100 ) , .A2( u1_u12_u7_n102 ) , .ZN( u1_u12_u7_n129 ) );
  NAND2_X1 u1_u12_u7_U64 (.A2( u1_u12_u7_n103 ) , .ZN( u1_u12_u7_n131 ) , .A1( u1_u12_u7_n95 ) );
  NAND2_X1 u1_u12_u7_U65 (.A1( u1_u12_u7_n100 ) , .ZN( u1_u12_u7_n138 ) , .A2( u1_u12_u7_n99 ) );
  NAND2_X1 u1_u12_u7_U66 (.ZN( u1_u12_u7_n132 ) , .A1( u1_u12_u7_n93 ) , .A2( u1_u12_u7_n96 ) );
  NAND2_X1 u1_u12_u7_U67 (.A1( u1_u12_u7_n100 ) , .ZN( u1_u12_u7_n148 ) , .A2( u1_u12_u7_n95 ) );
  NOR2_X1 u1_u12_u7_U68 (.A2( u1_u12_X_47 ) , .ZN( u1_u12_u7_n150 ) , .A1( u1_u12_u7_n163 ) );
  NOR2_X1 u1_u12_u7_U69 (.A2( u1_u12_X_43 ) , .A1( u1_u12_X_44 ) , .ZN( u1_u12_u7_n103 ) );
  AOI211_X1 u1_u12_u7_U7 (.ZN( u1_u12_u7_n116 ) , .A( u1_u12_u7_n155 ) , .C1( u1_u12_u7_n161 ) , .C2( u1_u12_u7_n171 ) , .B( u1_u12_u7_n94 ) );
  NOR2_X1 u1_u12_u7_U70 (.A2( u1_u12_X_48 ) , .A1( u1_u12_u7_n166 ) , .ZN( u1_u12_u7_n95 ) );
  NOR2_X1 u1_u12_u7_U71 (.A2( u1_u12_X_45 ) , .A1( u1_u12_X_48 ) , .ZN( u1_u12_u7_n99 ) );
  NOR2_X1 u1_u12_u7_U72 (.A2( u1_u12_X_44 ) , .A1( u1_u12_u7_n167 ) , .ZN( u1_u12_u7_n98 ) );
  NOR2_X1 u1_u12_u7_U73 (.A2( u1_u12_X_46 ) , .A1( u1_u12_X_47 ) , .ZN( u1_u12_u7_n152 ) );
  AND2_X1 u1_u12_u7_U74 (.A1( u1_u12_X_47 ) , .ZN( u1_u12_u7_n156 ) , .A2( u1_u12_u7_n163 ) );
  NAND2_X1 u1_u12_u7_U75 (.A2( u1_u12_X_46 ) , .A1( u1_u12_X_47 ) , .ZN( u1_u12_u7_n125 ) );
  AND2_X1 u1_u12_u7_U76 (.A2( u1_u12_X_45 ) , .A1( u1_u12_X_48 ) , .ZN( u1_u12_u7_n102 ) );
  AND2_X1 u1_u12_u7_U77 (.A2( u1_u12_X_43 ) , .A1( u1_u12_X_44 ) , .ZN( u1_u12_u7_n96 ) );
  AND2_X1 u1_u12_u7_U78 (.A1( u1_u12_X_44 ) , .ZN( u1_u12_u7_n100 ) , .A2( u1_u12_u7_n167 ) );
  AND2_X1 u1_u12_u7_U79 (.A1( u1_u12_X_48 ) , .A2( u1_u12_u7_n166 ) , .ZN( u1_u12_u7_n93 ) );
  OAI222_X1 u1_u12_u7_U8 (.C2( u1_u12_u7_n101 ) , .B2( u1_u12_u7_n111 ) , .A1( u1_u12_u7_n113 ) , .C1( u1_u12_u7_n146 ) , .A2( u1_u12_u7_n162 ) , .B1( u1_u12_u7_n164 ) , .ZN( u1_u12_u7_n94 ) );
  INV_X1 u1_u12_u7_U80 (.A( u1_u12_X_46 ) , .ZN( u1_u12_u7_n163 ) );
  INV_X1 u1_u12_u7_U81 (.A( u1_u12_X_43 ) , .ZN( u1_u12_u7_n167 ) );
  INV_X1 u1_u12_u7_U82 (.A( u1_u12_X_45 ) , .ZN( u1_u12_u7_n166 ) );
  NAND4_X1 u1_u12_u7_U83 (.ZN( u1_out12_5 ) , .A4( u1_u12_u7_n108 ) , .A3( u1_u12_u7_n109 ) , .A1( u1_u12_u7_n116 ) , .A2( u1_u12_u7_n123 ) );
  AOI22_X1 u1_u12_u7_U84 (.ZN( u1_u12_u7_n109 ) , .A2( u1_u12_u7_n126 ) , .B2( u1_u12_u7_n145 ) , .B1( u1_u12_u7_n156 ) , .A1( u1_u12_u7_n171 ) );
  NOR4_X1 u1_u12_u7_U85 (.A4( u1_u12_u7_n104 ) , .A3( u1_u12_u7_n105 ) , .A2( u1_u12_u7_n106 ) , .A1( u1_u12_u7_n107 ) , .ZN( u1_u12_u7_n108 ) );
  NAND4_X1 u1_u12_u7_U86 (.ZN( u1_out12_27 ) , .A4( u1_u12_u7_n118 ) , .A3( u1_u12_u7_n119 ) , .A2( u1_u12_u7_n120 ) , .A1( u1_u12_u7_n121 ) );
  OAI21_X1 u1_u12_u7_U87 (.ZN( u1_u12_u7_n121 ) , .B2( u1_u12_u7_n145 ) , .A( u1_u12_u7_n150 ) , .B1( u1_u12_u7_n174 ) );
  OAI21_X1 u1_u12_u7_U88 (.ZN( u1_u12_u7_n120 ) , .A( u1_u12_u7_n161 ) , .B2( u1_u12_u7_n170 ) , .B1( u1_u12_u7_n179 ) );
  NAND4_X1 u1_u12_u7_U89 (.ZN( u1_out12_21 ) , .A4( u1_u12_u7_n157 ) , .A3( u1_u12_u7_n158 ) , .A2( u1_u12_u7_n159 ) , .A1( u1_u12_u7_n160 ) );
  OAI221_X1 u1_u12_u7_U9 (.C1( u1_u12_u7_n101 ) , .C2( u1_u12_u7_n147 ) , .ZN( u1_u12_u7_n155 ) , .B2( u1_u12_u7_n162 ) , .A( u1_u12_u7_n91 ) , .B1( u1_u12_u7_n92 ) );
  OAI21_X1 u1_u12_u7_U90 (.B1( u1_u12_u7_n145 ) , .ZN( u1_u12_u7_n160 ) , .A( u1_u12_u7_n161 ) , .B2( u1_u12_u7_n177 ) );
  AOI22_X1 u1_u12_u7_U91 (.B2( u1_u12_u7_n149 ) , .B1( u1_u12_u7_n150 ) , .A2( u1_u12_u7_n151 ) , .A1( u1_u12_u7_n152 ) , .ZN( u1_u12_u7_n158 ) );
  NAND4_X1 u1_u12_u7_U92 (.ZN( u1_out12_15 ) , .A4( u1_u12_u7_n142 ) , .A3( u1_u12_u7_n143 ) , .A2( u1_u12_u7_n144 ) , .A1( u1_u12_u7_n178 ) );
  OR2_X1 u1_u12_u7_U93 (.A2( u1_u12_u7_n125 ) , .A1( u1_u12_u7_n129 ) , .ZN( u1_u12_u7_n144 ) );
  AOI22_X1 u1_u12_u7_U94 (.A2( u1_u12_u7_n126 ) , .ZN( u1_u12_u7_n143 ) , .B2( u1_u12_u7_n165 ) , .B1( u1_u12_u7_n173 ) , .A1( u1_u12_u7_n174 ) );
  NAND3_X1 u1_u12_u7_U95 (.A3( u1_u12_u7_n146 ) , .A2( u1_u12_u7_n147 ) , .A1( u1_u12_u7_n148 ) , .ZN( u1_u12_u7_n151 ) );
  NAND3_X1 u1_u12_u7_U96 (.A3( u1_u12_u7_n131 ) , .A2( u1_u12_u7_n132 ) , .A1( u1_u12_u7_n133 ) , .ZN( u1_u12_u7_n135 ) );
  XOR2_X1 u1_u13_U20 (.B( u1_K14_36 ) , .A( u1_R12_25 ) , .Z( u1_u13_X_36 ) );
  XOR2_X1 u1_u13_U21 (.B( u1_K14_35 ) , .A( u1_R12_24 ) , .Z( u1_u13_X_35 ) );
  XOR2_X1 u1_u13_U22 (.B( u1_K14_34 ) , .A( u1_R12_23 ) , .Z( u1_u13_X_34 ) );
  XOR2_X1 u1_u13_U23 (.B( u1_K14_33 ) , .A( u1_R12_22 ) , .Z( u1_u13_X_33 ) );
  XOR2_X1 u1_u13_U24 (.B( u1_K14_32 ) , .A( u1_R12_21 ) , .Z( u1_u13_X_32 ) );
  XOR2_X1 u1_u13_U25 (.B( u1_K14_31 ) , .A( u1_R12_20 ) , .Z( u1_u13_X_31 ) );
  XOR2_X1 u1_u13_U26 (.B( u1_K14_30 ) , .A( u1_R12_21 ) , .Z( u1_u13_X_30 ) );
  XOR2_X1 u1_u13_U28 (.B( u1_K14_29 ) , .A( u1_R12_20 ) , .Z( u1_u13_X_29 ) );
  XOR2_X1 u1_u13_U29 (.B( u1_K14_28 ) , .A( u1_R12_19 ) , .Z( u1_u13_X_28 ) );
  XOR2_X1 u1_u13_U30 (.B( u1_K14_27 ) , .A( u1_R12_18 ) , .Z( u1_u13_X_27 ) );
  XOR2_X1 u1_u13_U31 (.B( u1_K14_26 ) , .A( u1_R12_17 ) , .Z( u1_u13_X_26 ) );
  XOR2_X1 u1_u13_U32 (.B( u1_K14_25 ) , .A( u1_R12_16 ) , .Z( u1_u13_X_25 ) );
  OAI22_X1 u1_u13_u4_U10 (.B2( u1_u13_u4_n135 ) , .ZN( u1_u13_u4_n137 ) , .B1( u1_u13_u4_n153 ) , .A1( u1_u13_u4_n155 ) , .A2( u1_u13_u4_n171 ) );
  AND3_X1 u1_u13_u4_U11 (.A2( u1_u13_u4_n134 ) , .ZN( u1_u13_u4_n135 ) , .A3( u1_u13_u4_n145 ) , .A1( u1_u13_u4_n157 ) );
  NAND2_X1 u1_u13_u4_U12 (.ZN( u1_u13_u4_n132 ) , .A2( u1_u13_u4_n170 ) , .A1( u1_u13_u4_n173 ) );
  AOI21_X1 u1_u13_u4_U13 (.B2( u1_u13_u4_n160 ) , .B1( u1_u13_u4_n161 ) , .ZN( u1_u13_u4_n162 ) , .A( u1_u13_u4_n170 ) );
  AOI21_X1 u1_u13_u4_U14 (.ZN( u1_u13_u4_n107 ) , .B2( u1_u13_u4_n143 ) , .A( u1_u13_u4_n174 ) , .B1( u1_u13_u4_n184 ) );
  AOI21_X1 u1_u13_u4_U15 (.B2( u1_u13_u4_n158 ) , .B1( u1_u13_u4_n159 ) , .ZN( u1_u13_u4_n163 ) , .A( u1_u13_u4_n174 ) );
  AOI21_X1 u1_u13_u4_U16 (.A( u1_u13_u4_n153 ) , .B2( u1_u13_u4_n154 ) , .B1( u1_u13_u4_n155 ) , .ZN( u1_u13_u4_n165 ) );
  AOI21_X1 u1_u13_u4_U17 (.A( u1_u13_u4_n156 ) , .B2( u1_u13_u4_n157 ) , .ZN( u1_u13_u4_n164 ) , .B1( u1_u13_u4_n184 ) );
  INV_X1 u1_u13_u4_U18 (.A( u1_u13_u4_n138 ) , .ZN( u1_u13_u4_n170 ) );
  AND2_X1 u1_u13_u4_U19 (.A2( u1_u13_u4_n120 ) , .ZN( u1_u13_u4_n155 ) , .A1( u1_u13_u4_n160 ) );
  INV_X1 u1_u13_u4_U20 (.A( u1_u13_u4_n156 ) , .ZN( u1_u13_u4_n175 ) );
  NAND2_X1 u1_u13_u4_U21 (.A2( u1_u13_u4_n118 ) , .ZN( u1_u13_u4_n131 ) , .A1( u1_u13_u4_n147 ) );
  NAND2_X1 u1_u13_u4_U22 (.A1( u1_u13_u4_n119 ) , .A2( u1_u13_u4_n120 ) , .ZN( u1_u13_u4_n130 ) );
  NAND2_X1 u1_u13_u4_U23 (.ZN( u1_u13_u4_n117 ) , .A2( u1_u13_u4_n118 ) , .A1( u1_u13_u4_n148 ) );
  NAND2_X1 u1_u13_u4_U24 (.ZN( u1_u13_u4_n129 ) , .A1( u1_u13_u4_n134 ) , .A2( u1_u13_u4_n148 ) );
  AND3_X1 u1_u13_u4_U25 (.A1( u1_u13_u4_n119 ) , .A2( u1_u13_u4_n143 ) , .A3( u1_u13_u4_n154 ) , .ZN( u1_u13_u4_n161 ) );
  AND2_X1 u1_u13_u4_U26 (.A1( u1_u13_u4_n145 ) , .A2( u1_u13_u4_n147 ) , .ZN( u1_u13_u4_n159 ) );
  OR3_X1 u1_u13_u4_U27 (.A3( u1_u13_u4_n114 ) , .A2( u1_u13_u4_n115 ) , .A1( u1_u13_u4_n116 ) , .ZN( u1_u13_u4_n136 ) );
  AOI21_X1 u1_u13_u4_U28 (.A( u1_u13_u4_n113 ) , .ZN( u1_u13_u4_n116 ) , .B2( u1_u13_u4_n173 ) , .B1( u1_u13_u4_n174 ) );
  AOI21_X1 u1_u13_u4_U29 (.ZN( u1_u13_u4_n115 ) , .B2( u1_u13_u4_n145 ) , .B1( u1_u13_u4_n146 ) , .A( u1_u13_u4_n156 ) );
  NOR2_X1 u1_u13_u4_U3 (.ZN( u1_u13_u4_n121 ) , .A1( u1_u13_u4_n181 ) , .A2( u1_u13_u4_n182 ) );
  OAI22_X1 u1_u13_u4_U30 (.ZN( u1_u13_u4_n114 ) , .A2( u1_u13_u4_n121 ) , .B1( u1_u13_u4_n160 ) , .B2( u1_u13_u4_n170 ) , .A1( u1_u13_u4_n171 ) );
  INV_X1 u1_u13_u4_U31 (.A( u1_u13_u4_n158 ) , .ZN( u1_u13_u4_n182 ) );
  INV_X1 u1_u13_u4_U32 (.ZN( u1_u13_u4_n181 ) , .A( u1_u13_u4_n96 ) );
  INV_X1 u1_u13_u4_U33 (.A( u1_u13_u4_n144 ) , .ZN( u1_u13_u4_n179 ) );
  INV_X1 u1_u13_u4_U34 (.A( u1_u13_u4_n157 ) , .ZN( u1_u13_u4_n178 ) );
  NAND2_X1 u1_u13_u4_U35 (.A2( u1_u13_u4_n154 ) , .A1( u1_u13_u4_n96 ) , .ZN( u1_u13_u4_n97 ) );
  INV_X1 u1_u13_u4_U36 (.ZN( u1_u13_u4_n186 ) , .A( u1_u13_u4_n95 ) );
  OAI221_X1 u1_u13_u4_U37 (.C1( u1_u13_u4_n134 ) , .B1( u1_u13_u4_n158 ) , .B2( u1_u13_u4_n171 ) , .C2( u1_u13_u4_n173 ) , .A( u1_u13_u4_n94 ) , .ZN( u1_u13_u4_n95 ) );
  AOI222_X1 u1_u13_u4_U38 (.B2( u1_u13_u4_n132 ) , .A1( u1_u13_u4_n138 ) , .C2( u1_u13_u4_n175 ) , .A2( u1_u13_u4_n179 ) , .C1( u1_u13_u4_n181 ) , .B1( u1_u13_u4_n185 ) , .ZN( u1_u13_u4_n94 ) );
  INV_X1 u1_u13_u4_U39 (.A( u1_u13_u4_n113 ) , .ZN( u1_u13_u4_n185 ) );
  INV_X1 u1_u13_u4_U4 (.A( u1_u13_u4_n117 ) , .ZN( u1_u13_u4_n184 ) );
  INV_X1 u1_u13_u4_U40 (.A( u1_u13_u4_n143 ) , .ZN( u1_u13_u4_n183 ) );
  NOR2_X1 u1_u13_u4_U41 (.ZN( u1_u13_u4_n138 ) , .A1( u1_u13_u4_n168 ) , .A2( u1_u13_u4_n169 ) );
  NOR2_X1 u1_u13_u4_U42 (.A1( u1_u13_u4_n150 ) , .A2( u1_u13_u4_n152 ) , .ZN( u1_u13_u4_n153 ) );
  NOR2_X1 u1_u13_u4_U43 (.A2( u1_u13_u4_n128 ) , .A1( u1_u13_u4_n138 ) , .ZN( u1_u13_u4_n156 ) );
  AOI22_X1 u1_u13_u4_U44 (.B2( u1_u13_u4_n122 ) , .A1( u1_u13_u4_n123 ) , .ZN( u1_u13_u4_n124 ) , .B1( u1_u13_u4_n128 ) , .A2( u1_u13_u4_n172 ) );
  NAND2_X1 u1_u13_u4_U45 (.A2( u1_u13_u4_n120 ) , .ZN( u1_u13_u4_n123 ) , .A1( u1_u13_u4_n161 ) );
  INV_X1 u1_u13_u4_U46 (.A( u1_u13_u4_n153 ) , .ZN( u1_u13_u4_n172 ) );
  AOI22_X1 u1_u13_u4_U47 (.B2( u1_u13_u4_n132 ) , .A2( u1_u13_u4_n133 ) , .ZN( u1_u13_u4_n140 ) , .A1( u1_u13_u4_n150 ) , .B1( u1_u13_u4_n179 ) );
  NAND2_X1 u1_u13_u4_U48 (.ZN( u1_u13_u4_n133 ) , .A2( u1_u13_u4_n146 ) , .A1( u1_u13_u4_n154 ) );
  NAND2_X1 u1_u13_u4_U49 (.A1( u1_u13_u4_n103 ) , .ZN( u1_u13_u4_n154 ) , .A2( u1_u13_u4_n98 ) );
  NOR4_X1 u1_u13_u4_U5 (.A4( u1_u13_u4_n106 ) , .A3( u1_u13_u4_n107 ) , .A2( u1_u13_u4_n108 ) , .A1( u1_u13_u4_n109 ) , .ZN( u1_u13_u4_n110 ) );
  NAND2_X1 u1_u13_u4_U50 (.A1( u1_u13_u4_n101 ) , .ZN( u1_u13_u4_n158 ) , .A2( u1_u13_u4_n99 ) );
  AOI21_X1 u1_u13_u4_U51 (.ZN( u1_u13_u4_n127 ) , .A( u1_u13_u4_n136 ) , .B2( u1_u13_u4_n150 ) , .B1( u1_u13_u4_n180 ) );
  INV_X1 u1_u13_u4_U52 (.A( u1_u13_u4_n160 ) , .ZN( u1_u13_u4_n180 ) );
  NAND2_X1 u1_u13_u4_U53 (.A2( u1_u13_u4_n104 ) , .A1( u1_u13_u4_n105 ) , .ZN( u1_u13_u4_n146 ) );
  NAND2_X1 u1_u13_u4_U54 (.A2( u1_u13_u4_n101 ) , .A1( u1_u13_u4_n102 ) , .ZN( u1_u13_u4_n160 ) );
  NAND2_X1 u1_u13_u4_U55 (.ZN( u1_u13_u4_n134 ) , .A1( u1_u13_u4_n98 ) , .A2( u1_u13_u4_n99 ) );
  NAND2_X1 u1_u13_u4_U56 (.A1( u1_u13_u4_n103 ) , .A2( u1_u13_u4_n104 ) , .ZN( u1_u13_u4_n143 ) );
  NAND2_X1 u1_u13_u4_U57 (.A2( u1_u13_u4_n105 ) , .ZN( u1_u13_u4_n145 ) , .A1( u1_u13_u4_n98 ) );
  NAND2_X1 u1_u13_u4_U58 (.A1( u1_u13_u4_n100 ) , .A2( u1_u13_u4_n105 ) , .ZN( u1_u13_u4_n120 ) );
  NAND2_X1 u1_u13_u4_U59 (.A1( u1_u13_u4_n102 ) , .A2( u1_u13_u4_n104 ) , .ZN( u1_u13_u4_n148 ) );
  AOI21_X1 u1_u13_u4_U6 (.ZN( u1_u13_u4_n106 ) , .B2( u1_u13_u4_n146 ) , .B1( u1_u13_u4_n158 ) , .A( u1_u13_u4_n170 ) );
  NAND2_X1 u1_u13_u4_U60 (.A2( u1_u13_u4_n100 ) , .A1( u1_u13_u4_n103 ) , .ZN( u1_u13_u4_n157 ) );
  INV_X1 u1_u13_u4_U61 (.A( u1_u13_u4_n150 ) , .ZN( u1_u13_u4_n173 ) );
  INV_X1 u1_u13_u4_U62 (.A( u1_u13_u4_n152 ) , .ZN( u1_u13_u4_n171 ) );
  NAND2_X1 u1_u13_u4_U63 (.A1( u1_u13_u4_n100 ) , .ZN( u1_u13_u4_n118 ) , .A2( u1_u13_u4_n99 ) );
  NAND2_X1 u1_u13_u4_U64 (.A2( u1_u13_u4_n100 ) , .A1( u1_u13_u4_n102 ) , .ZN( u1_u13_u4_n144 ) );
  NAND2_X1 u1_u13_u4_U65 (.A2( u1_u13_u4_n101 ) , .A1( u1_u13_u4_n105 ) , .ZN( u1_u13_u4_n96 ) );
  INV_X1 u1_u13_u4_U66 (.A( u1_u13_u4_n128 ) , .ZN( u1_u13_u4_n174 ) );
  NAND2_X1 u1_u13_u4_U67 (.A2( u1_u13_u4_n102 ) , .ZN( u1_u13_u4_n119 ) , .A1( u1_u13_u4_n98 ) );
  NAND2_X1 u1_u13_u4_U68 (.A2( u1_u13_u4_n101 ) , .A1( u1_u13_u4_n103 ) , .ZN( u1_u13_u4_n147 ) );
  NAND2_X1 u1_u13_u4_U69 (.A2( u1_u13_u4_n104 ) , .ZN( u1_u13_u4_n113 ) , .A1( u1_u13_u4_n99 ) );
  AOI21_X1 u1_u13_u4_U7 (.ZN( u1_u13_u4_n108 ) , .B2( u1_u13_u4_n134 ) , .B1( u1_u13_u4_n155 ) , .A( u1_u13_u4_n156 ) );
  NOR2_X1 u1_u13_u4_U70 (.A2( u1_u13_X_28 ) , .ZN( u1_u13_u4_n150 ) , .A1( u1_u13_u4_n168 ) );
  NOR2_X1 u1_u13_u4_U71 (.A2( u1_u13_X_29 ) , .ZN( u1_u13_u4_n152 ) , .A1( u1_u13_u4_n169 ) );
  NOR2_X1 u1_u13_u4_U72 (.A2( u1_u13_X_30 ) , .ZN( u1_u13_u4_n105 ) , .A1( u1_u13_u4_n176 ) );
  NOR2_X1 u1_u13_u4_U73 (.A2( u1_u13_X_26 ) , .ZN( u1_u13_u4_n100 ) , .A1( u1_u13_u4_n177 ) );
  NOR2_X1 u1_u13_u4_U74 (.A2( u1_u13_X_28 ) , .A1( u1_u13_X_29 ) , .ZN( u1_u13_u4_n128 ) );
  NOR2_X1 u1_u13_u4_U75 (.A2( u1_u13_X_27 ) , .A1( u1_u13_X_30 ) , .ZN( u1_u13_u4_n102 ) );
  NOR2_X1 u1_u13_u4_U76 (.A2( u1_u13_X_25 ) , .A1( u1_u13_X_26 ) , .ZN( u1_u13_u4_n98 ) );
  AND2_X1 u1_u13_u4_U77 (.A2( u1_u13_X_25 ) , .A1( u1_u13_X_26 ) , .ZN( u1_u13_u4_n104 ) );
  AND2_X1 u1_u13_u4_U78 (.A1( u1_u13_X_30 ) , .A2( u1_u13_u4_n176 ) , .ZN( u1_u13_u4_n99 ) );
  AND2_X1 u1_u13_u4_U79 (.A1( u1_u13_X_26 ) , .ZN( u1_u13_u4_n101 ) , .A2( u1_u13_u4_n177 ) );
  AOI21_X1 u1_u13_u4_U8 (.ZN( u1_u13_u4_n109 ) , .A( u1_u13_u4_n153 ) , .B1( u1_u13_u4_n159 ) , .B2( u1_u13_u4_n184 ) );
  AND2_X1 u1_u13_u4_U80 (.A1( u1_u13_X_27 ) , .A2( u1_u13_X_30 ) , .ZN( u1_u13_u4_n103 ) );
  INV_X1 u1_u13_u4_U81 (.A( u1_u13_X_28 ) , .ZN( u1_u13_u4_n169 ) );
  INV_X1 u1_u13_u4_U82 (.A( u1_u13_X_29 ) , .ZN( u1_u13_u4_n168 ) );
  INV_X1 u1_u13_u4_U83 (.A( u1_u13_X_25 ) , .ZN( u1_u13_u4_n177 ) );
  INV_X1 u1_u13_u4_U84 (.A( u1_u13_X_27 ) , .ZN( u1_u13_u4_n176 ) );
  NAND4_X1 u1_u13_u4_U85 (.ZN( u1_out13_25 ) , .A4( u1_u13_u4_n139 ) , .A3( u1_u13_u4_n140 ) , .A2( u1_u13_u4_n141 ) , .A1( u1_u13_u4_n142 ) );
  OAI21_X1 u1_u13_u4_U86 (.A( u1_u13_u4_n128 ) , .B2( u1_u13_u4_n129 ) , .B1( u1_u13_u4_n130 ) , .ZN( u1_u13_u4_n142 ) );
  OAI21_X1 u1_u13_u4_U87 (.B2( u1_u13_u4_n131 ) , .ZN( u1_u13_u4_n141 ) , .A( u1_u13_u4_n175 ) , .B1( u1_u13_u4_n183 ) );
  NAND4_X1 u1_u13_u4_U88 (.ZN( u1_out13_14 ) , .A4( u1_u13_u4_n124 ) , .A3( u1_u13_u4_n125 ) , .A2( u1_u13_u4_n126 ) , .A1( u1_u13_u4_n127 ) );
  AOI22_X1 u1_u13_u4_U89 (.B2( u1_u13_u4_n117 ) , .ZN( u1_u13_u4_n126 ) , .A1( u1_u13_u4_n129 ) , .B1( u1_u13_u4_n152 ) , .A2( u1_u13_u4_n175 ) );
  AOI211_X1 u1_u13_u4_U9 (.B( u1_u13_u4_n136 ) , .A( u1_u13_u4_n137 ) , .C2( u1_u13_u4_n138 ) , .ZN( u1_u13_u4_n139 ) , .C1( u1_u13_u4_n182 ) );
  AOI22_X1 u1_u13_u4_U90 (.ZN( u1_u13_u4_n125 ) , .B2( u1_u13_u4_n131 ) , .A2( u1_u13_u4_n132 ) , .B1( u1_u13_u4_n138 ) , .A1( u1_u13_u4_n178 ) );
  NAND4_X1 u1_u13_u4_U91 (.ZN( u1_out13_8 ) , .A4( u1_u13_u4_n110 ) , .A3( u1_u13_u4_n111 ) , .A2( u1_u13_u4_n112 ) , .A1( u1_u13_u4_n186 ) );
  NAND2_X1 u1_u13_u4_U92 (.ZN( u1_u13_u4_n112 ) , .A2( u1_u13_u4_n130 ) , .A1( u1_u13_u4_n150 ) );
  AOI22_X1 u1_u13_u4_U93 (.ZN( u1_u13_u4_n111 ) , .B2( u1_u13_u4_n132 ) , .A1( u1_u13_u4_n152 ) , .B1( u1_u13_u4_n178 ) , .A2( u1_u13_u4_n97 ) );
  AOI22_X1 u1_u13_u4_U94 (.B2( u1_u13_u4_n149 ) , .B1( u1_u13_u4_n150 ) , .A2( u1_u13_u4_n151 ) , .A1( u1_u13_u4_n152 ) , .ZN( u1_u13_u4_n167 ) );
  NOR4_X1 u1_u13_u4_U95 (.A4( u1_u13_u4_n162 ) , .A3( u1_u13_u4_n163 ) , .A2( u1_u13_u4_n164 ) , .A1( u1_u13_u4_n165 ) , .ZN( u1_u13_u4_n166 ) );
  NAND3_X1 u1_u13_u4_U96 (.ZN( u1_out13_3 ) , .A3( u1_u13_u4_n166 ) , .A1( u1_u13_u4_n167 ) , .A2( u1_u13_u4_n186 ) );
  NAND3_X1 u1_u13_u4_U97 (.A3( u1_u13_u4_n146 ) , .A2( u1_u13_u4_n147 ) , .A1( u1_u13_u4_n148 ) , .ZN( u1_u13_u4_n149 ) );
  NAND3_X1 u1_u13_u4_U98 (.A3( u1_u13_u4_n143 ) , .A2( u1_u13_u4_n144 ) , .A1( u1_u13_u4_n145 ) , .ZN( u1_u13_u4_n151 ) );
  NAND3_X1 u1_u13_u4_U99 (.A3( u1_u13_u4_n121 ) , .ZN( u1_u13_u4_n122 ) , .A2( u1_u13_u4_n144 ) , .A1( u1_u13_u4_n154 ) );
  INV_X1 u1_u13_u5_U10 (.A( u1_u13_u5_n121 ) , .ZN( u1_u13_u5_n177 ) );
  AOI222_X1 u1_u13_u5_U100 (.ZN( u1_u13_u5_n113 ) , .A1( u1_u13_u5_n131 ) , .C1( u1_u13_u5_n148 ) , .B2( u1_u13_u5_n174 ) , .C2( u1_u13_u5_n178 ) , .A2( u1_u13_u5_n179 ) , .B1( u1_u13_u5_n99 ) );
  NAND4_X1 u1_u13_u5_U101 (.ZN( u1_out13_11 ) , .A4( u1_u13_u5_n143 ) , .A3( u1_u13_u5_n144 ) , .A2( u1_u13_u5_n169 ) , .A1( u1_u13_u5_n196 ) );
  AOI22_X1 u1_u13_u5_U102 (.A2( u1_u13_u5_n132 ) , .ZN( u1_u13_u5_n144 ) , .B2( u1_u13_u5_n145 ) , .B1( u1_u13_u5_n184 ) , .A1( u1_u13_u5_n194 ) );
  NOR3_X1 u1_u13_u5_U103 (.A3( u1_u13_u5_n141 ) , .A1( u1_u13_u5_n142 ) , .ZN( u1_u13_u5_n143 ) , .A2( u1_u13_u5_n191 ) );
  NAND3_X1 u1_u13_u5_U104 (.A2( u1_u13_u5_n154 ) , .A3( u1_u13_u5_n158 ) , .A1( u1_u13_u5_n161 ) , .ZN( u1_u13_u5_n99 ) );
  NOR2_X1 u1_u13_u5_U11 (.ZN( u1_u13_u5_n160 ) , .A2( u1_u13_u5_n173 ) , .A1( u1_u13_u5_n177 ) );
  INV_X1 u1_u13_u5_U12 (.A( u1_u13_u5_n150 ) , .ZN( u1_u13_u5_n174 ) );
  AOI21_X1 u1_u13_u5_U13 (.A( u1_u13_u5_n160 ) , .B2( u1_u13_u5_n161 ) , .ZN( u1_u13_u5_n162 ) , .B1( u1_u13_u5_n192 ) );
  INV_X1 u1_u13_u5_U14 (.A( u1_u13_u5_n159 ) , .ZN( u1_u13_u5_n192 ) );
  AOI21_X1 u1_u13_u5_U15 (.A( u1_u13_u5_n156 ) , .B2( u1_u13_u5_n157 ) , .B1( u1_u13_u5_n158 ) , .ZN( u1_u13_u5_n163 ) );
  AOI21_X1 u1_u13_u5_U16 (.B2( u1_u13_u5_n139 ) , .B1( u1_u13_u5_n140 ) , .ZN( u1_u13_u5_n141 ) , .A( u1_u13_u5_n150 ) );
  OAI21_X1 u1_u13_u5_U17 (.A( u1_u13_u5_n133 ) , .B2( u1_u13_u5_n134 ) , .B1( u1_u13_u5_n135 ) , .ZN( u1_u13_u5_n142 ) );
  OAI21_X1 u1_u13_u5_U18 (.ZN( u1_u13_u5_n133 ) , .B2( u1_u13_u5_n147 ) , .A( u1_u13_u5_n173 ) , .B1( u1_u13_u5_n188 ) );
  NAND2_X1 u1_u13_u5_U19 (.A2( u1_u13_u5_n119 ) , .A1( u1_u13_u5_n123 ) , .ZN( u1_u13_u5_n137 ) );
  INV_X1 u1_u13_u5_U20 (.A( u1_u13_u5_n155 ) , .ZN( u1_u13_u5_n194 ) );
  NAND2_X1 u1_u13_u5_U21 (.A1( u1_u13_u5_n121 ) , .ZN( u1_u13_u5_n132 ) , .A2( u1_u13_u5_n172 ) );
  NAND2_X1 u1_u13_u5_U22 (.A2( u1_u13_u5_n122 ) , .ZN( u1_u13_u5_n136 ) , .A1( u1_u13_u5_n154 ) );
  NAND2_X1 u1_u13_u5_U23 (.A2( u1_u13_u5_n119 ) , .A1( u1_u13_u5_n120 ) , .ZN( u1_u13_u5_n159 ) );
  INV_X1 u1_u13_u5_U24 (.A( u1_u13_u5_n156 ) , .ZN( u1_u13_u5_n175 ) );
  INV_X1 u1_u13_u5_U25 (.A( u1_u13_u5_n158 ) , .ZN( u1_u13_u5_n188 ) );
  INV_X1 u1_u13_u5_U26 (.A( u1_u13_u5_n152 ) , .ZN( u1_u13_u5_n179 ) );
  INV_X1 u1_u13_u5_U27 (.A( u1_u13_u5_n140 ) , .ZN( u1_u13_u5_n182 ) );
  INV_X1 u1_u13_u5_U28 (.A( u1_u13_u5_n151 ) , .ZN( u1_u13_u5_n183 ) );
  INV_X1 u1_u13_u5_U29 (.A( u1_u13_u5_n123 ) , .ZN( u1_u13_u5_n185 ) );
  NOR2_X1 u1_u13_u5_U3 (.ZN( u1_u13_u5_n134 ) , .A1( u1_u13_u5_n183 ) , .A2( u1_u13_u5_n190 ) );
  INV_X1 u1_u13_u5_U30 (.A( u1_u13_u5_n161 ) , .ZN( u1_u13_u5_n184 ) );
  INV_X1 u1_u13_u5_U31 (.A( u1_u13_u5_n139 ) , .ZN( u1_u13_u5_n189 ) );
  INV_X1 u1_u13_u5_U32 (.A( u1_u13_u5_n157 ) , .ZN( u1_u13_u5_n190 ) );
  INV_X1 u1_u13_u5_U33 (.A( u1_u13_u5_n120 ) , .ZN( u1_u13_u5_n193 ) );
  NAND2_X1 u1_u13_u5_U34 (.ZN( u1_u13_u5_n111 ) , .A1( u1_u13_u5_n140 ) , .A2( u1_u13_u5_n155 ) );
  INV_X1 u1_u13_u5_U35 (.A( u1_u13_u5_n117 ) , .ZN( u1_u13_u5_n196 ) );
  OAI221_X1 u1_u13_u5_U36 (.A( u1_u13_u5_n116 ) , .ZN( u1_u13_u5_n117 ) , .B2( u1_u13_u5_n119 ) , .C1( u1_u13_u5_n153 ) , .C2( u1_u13_u5_n158 ) , .B1( u1_u13_u5_n172 ) );
  AOI222_X1 u1_u13_u5_U37 (.ZN( u1_u13_u5_n116 ) , .B2( u1_u13_u5_n145 ) , .C1( u1_u13_u5_n148 ) , .A2( u1_u13_u5_n174 ) , .C2( u1_u13_u5_n177 ) , .B1( u1_u13_u5_n187 ) , .A1( u1_u13_u5_n193 ) );
  INV_X1 u1_u13_u5_U38 (.A( u1_u13_u5_n115 ) , .ZN( u1_u13_u5_n187 ) );
  NOR2_X1 u1_u13_u5_U39 (.ZN( u1_u13_u5_n100 ) , .A1( u1_u13_u5_n170 ) , .A2( u1_u13_u5_n180 ) );
  INV_X1 u1_u13_u5_U4 (.A( u1_u13_u5_n138 ) , .ZN( u1_u13_u5_n191 ) );
  AOI22_X1 u1_u13_u5_U40 (.B2( u1_u13_u5_n131 ) , .A2( u1_u13_u5_n146 ) , .ZN( u1_u13_u5_n169 ) , .B1( u1_u13_u5_n174 ) , .A1( u1_u13_u5_n185 ) );
  NOR2_X1 u1_u13_u5_U41 (.A1( u1_u13_u5_n146 ) , .ZN( u1_u13_u5_n150 ) , .A2( u1_u13_u5_n173 ) );
  AOI21_X1 u1_u13_u5_U42 (.A( u1_u13_u5_n118 ) , .B2( u1_u13_u5_n145 ) , .ZN( u1_u13_u5_n168 ) , .B1( u1_u13_u5_n186 ) );
  INV_X1 u1_u13_u5_U43 (.A( u1_u13_u5_n122 ) , .ZN( u1_u13_u5_n186 ) );
  NOR2_X1 u1_u13_u5_U44 (.A1( u1_u13_u5_n146 ) , .ZN( u1_u13_u5_n152 ) , .A2( u1_u13_u5_n176 ) );
  NOR2_X1 u1_u13_u5_U45 (.A1( u1_u13_u5_n115 ) , .ZN( u1_u13_u5_n118 ) , .A2( u1_u13_u5_n153 ) );
  NOR2_X1 u1_u13_u5_U46 (.A2( u1_u13_u5_n145 ) , .ZN( u1_u13_u5_n156 ) , .A1( u1_u13_u5_n174 ) );
  NOR2_X1 u1_u13_u5_U47 (.ZN( u1_u13_u5_n121 ) , .A2( u1_u13_u5_n145 ) , .A1( u1_u13_u5_n176 ) );
  AOI22_X1 u1_u13_u5_U48 (.ZN( u1_u13_u5_n114 ) , .A2( u1_u13_u5_n137 ) , .A1( u1_u13_u5_n145 ) , .B2( u1_u13_u5_n175 ) , .B1( u1_u13_u5_n193 ) );
  OAI211_X1 u1_u13_u5_U49 (.B( u1_u13_u5_n124 ) , .A( u1_u13_u5_n125 ) , .C2( u1_u13_u5_n126 ) , .C1( u1_u13_u5_n127 ) , .ZN( u1_u13_u5_n128 ) );
  OAI21_X1 u1_u13_u5_U5 (.B2( u1_u13_u5_n136 ) , .B1( u1_u13_u5_n137 ) , .ZN( u1_u13_u5_n138 ) , .A( u1_u13_u5_n177 ) );
  NOR3_X1 u1_u13_u5_U50 (.ZN( u1_u13_u5_n127 ) , .A1( u1_u13_u5_n136 ) , .A3( u1_u13_u5_n148 ) , .A2( u1_u13_u5_n182 ) );
  OAI21_X1 u1_u13_u5_U51 (.ZN( u1_u13_u5_n124 ) , .A( u1_u13_u5_n177 ) , .B2( u1_u13_u5_n183 ) , .B1( u1_u13_u5_n189 ) );
  OAI21_X1 u1_u13_u5_U52 (.ZN( u1_u13_u5_n125 ) , .A( u1_u13_u5_n174 ) , .B2( u1_u13_u5_n185 ) , .B1( u1_u13_u5_n190 ) );
  AOI21_X1 u1_u13_u5_U53 (.A( u1_u13_u5_n153 ) , .B2( u1_u13_u5_n154 ) , .B1( u1_u13_u5_n155 ) , .ZN( u1_u13_u5_n164 ) );
  AOI21_X1 u1_u13_u5_U54 (.ZN( u1_u13_u5_n110 ) , .B1( u1_u13_u5_n122 ) , .B2( u1_u13_u5_n139 ) , .A( u1_u13_u5_n153 ) );
  INV_X1 u1_u13_u5_U55 (.A( u1_u13_u5_n153 ) , .ZN( u1_u13_u5_n176 ) );
  INV_X1 u1_u13_u5_U56 (.A( u1_u13_u5_n126 ) , .ZN( u1_u13_u5_n173 ) );
  AND2_X1 u1_u13_u5_U57 (.A2( u1_u13_u5_n104 ) , .A1( u1_u13_u5_n107 ) , .ZN( u1_u13_u5_n147 ) );
  AND2_X1 u1_u13_u5_U58 (.A2( u1_u13_u5_n104 ) , .A1( u1_u13_u5_n108 ) , .ZN( u1_u13_u5_n148 ) );
  NAND2_X1 u1_u13_u5_U59 (.A1( u1_u13_u5_n105 ) , .A2( u1_u13_u5_n106 ) , .ZN( u1_u13_u5_n158 ) );
  INV_X1 u1_u13_u5_U6 (.A( u1_u13_u5_n135 ) , .ZN( u1_u13_u5_n178 ) );
  NAND2_X1 u1_u13_u5_U60 (.A2( u1_u13_u5_n108 ) , .A1( u1_u13_u5_n109 ) , .ZN( u1_u13_u5_n139 ) );
  NAND2_X1 u1_u13_u5_U61 (.A1( u1_u13_u5_n106 ) , .A2( u1_u13_u5_n108 ) , .ZN( u1_u13_u5_n119 ) );
  NAND2_X1 u1_u13_u5_U62 (.A2( u1_u13_u5_n103 ) , .A1( u1_u13_u5_n105 ) , .ZN( u1_u13_u5_n140 ) );
  NAND2_X1 u1_u13_u5_U63 (.A2( u1_u13_u5_n104 ) , .A1( u1_u13_u5_n105 ) , .ZN( u1_u13_u5_n155 ) );
  NAND2_X1 u1_u13_u5_U64 (.A2( u1_u13_u5_n106 ) , .A1( u1_u13_u5_n107 ) , .ZN( u1_u13_u5_n122 ) );
  NAND2_X1 u1_u13_u5_U65 (.A2( u1_u13_u5_n100 ) , .A1( u1_u13_u5_n106 ) , .ZN( u1_u13_u5_n115 ) );
  NAND2_X1 u1_u13_u5_U66 (.A2( u1_u13_u5_n100 ) , .A1( u1_u13_u5_n103 ) , .ZN( u1_u13_u5_n161 ) );
  NAND2_X1 u1_u13_u5_U67 (.A1( u1_u13_u5_n105 ) , .A2( u1_u13_u5_n109 ) , .ZN( u1_u13_u5_n154 ) );
  INV_X1 u1_u13_u5_U68 (.A( u1_u13_u5_n146 ) , .ZN( u1_u13_u5_n172 ) );
  NAND2_X1 u1_u13_u5_U69 (.A1( u1_u13_u5_n103 ) , .A2( u1_u13_u5_n108 ) , .ZN( u1_u13_u5_n123 ) );
  OAI22_X1 u1_u13_u5_U7 (.B2( u1_u13_u5_n149 ) , .B1( u1_u13_u5_n150 ) , .A2( u1_u13_u5_n151 ) , .A1( u1_u13_u5_n152 ) , .ZN( u1_u13_u5_n165 ) );
  NAND2_X1 u1_u13_u5_U70 (.A2( u1_u13_u5_n103 ) , .A1( u1_u13_u5_n107 ) , .ZN( u1_u13_u5_n151 ) );
  NAND2_X1 u1_u13_u5_U71 (.A2( u1_u13_u5_n107 ) , .A1( u1_u13_u5_n109 ) , .ZN( u1_u13_u5_n120 ) );
  NAND2_X1 u1_u13_u5_U72 (.A2( u1_u13_u5_n100 ) , .A1( u1_u13_u5_n109 ) , .ZN( u1_u13_u5_n157 ) );
  AND2_X1 u1_u13_u5_U73 (.A2( u1_u13_u5_n100 ) , .A1( u1_u13_u5_n104 ) , .ZN( u1_u13_u5_n131 ) );
  INV_X1 u1_u13_u5_U74 (.A( u1_u13_u5_n102 ) , .ZN( u1_u13_u5_n195 ) );
  OAI221_X1 u1_u13_u5_U75 (.A( u1_u13_u5_n101 ) , .ZN( u1_u13_u5_n102 ) , .C2( u1_u13_u5_n115 ) , .C1( u1_u13_u5_n126 ) , .B1( u1_u13_u5_n134 ) , .B2( u1_u13_u5_n160 ) );
  OAI21_X1 u1_u13_u5_U76 (.ZN( u1_u13_u5_n101 ) , .B1( u1_u13_u5_n137 ) , .A( u1_u13_u5_n146 ) , .B2( u1_u13_u5_n147 ) );
  NOR2_X1 u1_u13_u5_U77 (.A2( u1_u13_X_34 ) , .A1( u1_u13_X_35 ) , .ZN( u1_u13_u5_n145 ) );
  NOR2_X1 u1_u13_u5_U78 (.A2( u1_u13_X_34 ) , .ZN( u1_u13_u5_n146 ) , .A1( u1_u13_u5_n171 ) );
  NOR2_X1 u1_u13_u5_U79 (.A2( u1_u13_X_31 ) , .A1( u1_u13_X_32 ) , .ZN( u1_u13_u5_n103 ) );
  NOR3_X1 u1_u13_u5_U8 (.A2( u1_u13_u5_n147 ) , .A1( u1_u13_u5_n148 ) , .ZN( u1_u13_u5_n149 ) , .A3( u1_u13_u5_n194 ) );
  NOR2_X1 u1_u13_u5_U80 (.A2( u1_u13_X_36 ) , .ZN( u1_u13_u5_n105 ) , .A1( u1_u13_u5_n180 ) );
  NOR2_X1 u1_u13_u5_U81 (.A2( u1_u13_X_33 ) , .ZN( u1_u13_u5_n108 ) , .A1( u1_u13_u5_n170 ) );
  NOR2_X1 u1_u13_u5_U82 (.A2( u1_u13_X_33 ) , .A1( u1_u13_X_36 ) , .ZN( u1_u13_u5_n107 ) );
  NOR2_X1 u1_u13_u5_U83 (.A2( u1_u13_X_31 ) , .ZN( u1_u13_u5_n104 ) , .A1( u1_u13_u5_n181 ) );
  NAND2_X1 u1_u13_u5_U84 (.A2( u1_u13_X_34 ) , .A1( u1_u13_X_35 ) , .ZN( u1_u13_u5_n153 ) );
  NAND2_X1 u1_u13_u5_U85 (.A1( u1_u13_X_34 ) , .ZN( u1_u13_u5_n126 ) , .A2( u1_u13_u5_n171 ) );
  AND2_X1 u1_u13_u5_U86 (.A1( u1_u13_X_31 ) , .A2( u1_u13_X_32 ) , .ZN( u1_u13_u5_n106 ) );
  AND2_X1 u1_u13_u5_U87 (.A1( u1_u13_X_31 ) , .ZN( u1_u13_u5_n109 ) , .A2( u1_u13_u5_n181 ) );
  INV_X1 u1_u13_u5_U88 (.A( u1_u13_X_33 ) , .ZN( u1_u13_u5_n180 ) );
  INV_X1 u1_u13_u5_U89 (.A( u1_u13_X_35 ) , .ZN( u1_u13_u5_n171 ) );
  NOR2_X1 u1_u13_u5_U9 (.ZN( u1_u13_u5_n135 ) , .A1( u1_u13_u5_n173 ) , .A2( u1_u13_u5_n176 ) );
  INV_X1 u1_u13_u5_U90 (.A( u1_u13_X_36 ) , .ZN( u1_u13_u5_n170 ) );
  INV_X1 u1_u13_u5_U91 (.A( u1_u13_X_32 ) , .ZN( u1_u13_u5_n181 ) );
  NAND4_X1 u1_u13_u5_U92 (.ZN( u1_out13_29 ) , .A4( u1_u13_u5_n129 ) , .A3( u1_u13_u5_n130 ) , .A2( u1_u13_u5_n168 ) , .A1( u1_u13_u5_n196 ) );
  AOI221_X1 u1_u13_u5_U93 (.A( u1_u13_u5_n128 ) , .ZN( u1_u13_u5_n129 ) , .C2( u1_u13_u5_n132 ) , .B2( u1_u13_u5_n159 ) , .B1( u1_u13_u5_n176 ) , .C1( u1_u13_u5_n184 ) );
  AOI222_X1 u1_u13_u5_U94 (.ZN( u1_u13_u5_n130 ) , .A2( u1_u13_u5_n146 ) , .B1( u1_u13_u5_n147 ) , .C2( u1_u13_u5_n175 ) , .B2( u1_u13_u5_n179 ) , .A1( u1_u13_u5_n188 ) , .C1( u1_u13_u5_n194 ) );
  NAND4_X1 u1_u13_u5_U95 (.ZN( u1_out13_19 ) , .A4( u1_u13_u5_n166 ) , .A3( u1_u13_u5_n167 ) , .A2( u1_u13_u5_n168 ) , .A1( u1_u13_u5_n169 ) );
  AOI22_X1 u1_u13_u5_U96 (.B2( u1_u13_u5_n145 ) , .A2( u1_u13_u5_n146 ) , .ZN( u1_u13_u5_n167 ) , .B1( u1_u13_u5_n182 ) , .A1( u1_u13_u5_n189 ) );
  NOR4_X1 u1_u13_u5_U97 (.A4( u1_u13_u5_n162 ) , .A3( u1_u13_u5_n163 ) , .A2( u1_u13_u5_n164 ) , .A1( u1_u13_u5_n165 ) , .ZN( u1_u13_u5_n166 ) );
  NAND4_X1 u1_u13_u5_U98 (.ZN( u1_out13_4 ) , .A4( u1_u13_u5_n112 ) , .A2( u1_u13_u5_n113 ) , .A1( u1_u13_u5_n114 ) , .A3( u1_u13_u5_n195 ) );
  AOI211_X1 u1_u13_u5_U99 (.A( u1_u13_u5_n110 ) , .C1( u1_u13_u5_n111 ) , .ZN( u1_u13_u5_n112 ) , .B( u1_u13_u5_n118 ) , .C2( u1_u13_u5_n177 ) );
  XOR2_X1 u1_u1_U13 (.B( u1_K2_42 ) , .A( u1_R0_29 ) , .Z( u1_u1_X_42 ) );
  XOR2_X1 u1_u1_U14 (.B( u1_K2_41 ) , .A( u1_R0_28 ) , .Z( u1_u1_X_41 ) );
  XOR2_X1 u1_u1_U15 (.B( u1_K2_40 ) , .A( u1_R0_27 ) , .Z( u1_u1_X_40 ) );
  XOR2_X1 u1_u1_U17 (.B( u1_K2_39 ) , .A( u1_R0_26 ) , .Z( u1_u1_X_39 ) );
  XOR2_X1 u1_u1_U18 (.B( u1_K2_38 ) , .A( u1_R0_25 ) , .Z( u1_u1_X_38 ) );
  XOR2_X1 u1_u1_U19 (.B( u1_K2_37 ) , .A( u1_R0_24 ) , .Z( u1_u1_X_37 ) );
  XOR2_X1 u1_u1_U26 (.B( u1_K2_30 ) , .A( u1_R0_21 ) , .Z( u1_u1_X_30 ) );
  XOR2_X1 u1_u1_U28 (.B( u1_K2_29 ) , .A( u1_R0_20 ) , .Z( u1_u1_X_29 ) );
  XOR2_X1 u1_u1_U29 (.B( u1_K2_28 ) , .A( u1_R0_19 ) , .Z( u1_u1_X_28 ) );
  XOR2_X1 u1_u1_U30 (.B( u1_K2_27 ) , .A( u1_R0_18 ) , .Z( u1_u1_X_27 ) );
  XOR2_X1 u1_u1_U31 (.B( u1_K2_26 ) , .A( u1_R0_17 ) , .Z( u1_u1_X_26 ) );
  XOR2_X1 u1_u1_U32 (.B( u1_K2_25 ) , .A( u1_R0_16 ) , .Z( u1_u1_X_25 ) );
  OAI22_X1 u1_u1_u4_U10 (.B2( u1_u1_u4_n135 ) , .ZN( u1_u1_u4_n137 ) , .B1( u1_u1_u4_n153 ) , .A1( u1_u1_u4_n155 ) , .A2( u1_u1_u4_n171 ) );
  AND3_X1 u1_u1_u4_U11 (.A2( u1_u1_u4_n134 ) , .ZN( u1_u1_u4_n135 ) , .A3( u1_u1_u4_n145 ) , .A1( u1_u1_u4_n157 ) );
  NAND2_X1 u1_u1_u4_U12 (.ZN( u1_u1_u4_n132 ) , .A2( u1_u1_u4_n170 ) , .A1( u1_u1_u4_n173 ) );
  AOI21_X1 u1_u1_u4_U13 (.B2( u1_u1_u4_n160 ) , .B1( u1_u1_u4_n161 ) , .ZN( u1_u1_u4_n162 ) , .A( u1_u1_u4_n170 ) );
  AOI21_X1 u1_u1_u4_U14 (.ZN( u1_u1_u4_n107 ) , .B2( u1_u1_u4_n143 ) , .A( u1_u1_u4_n174 ) , .B1( u1_u1_u4_n184 ) );
  AOI21_X1 u1_u1_u4_U15 (.B2( u1_u1_u4_n158 ) , .B1( u1_u1_u4_n159 ) , .ZN( u1_u1_u4_n163 ) , .A( u1_u1_u4_n174 ) );
  AOI21_X1 u1_u1_u4_U16 (.A( u1_u1_u4_n153 ) , .B2( u1_u1_u4_n154 ) , .B1( u1_u1_u4_n155 ) , .ZN( u1_u1_u4_n165 ) );
  AOI21_X1 u1_u1_u4_U17 (.A( u1_u1_u4_n156 ) , .B2( u1_u1_u4_n157 ) , .ZN( u1_u1_u4_n164 ) , .B1( u1_u1_u4_n184 ) );
  INV_X1 u1_u1_u4_U18 (.A( u1_u1_u4_n138 ) , .ZN( u1_u1_u4_n170 ) );
  AND2_X1 u1_u1_u4_U19 (.A2( u1_u1_u4_n120 ) , .ZN( u1_u1_u4_n155 ) , .A1( u1_u1_u4_n160 ) );
  INV_X1 u1_u1_u4_U20 (.A( u1_u1_u4_n156 ) , .ZN( u1_u1_u4_n175 ) );
  NAND2_X1 u1_u1_u4_U21 (.A2( u1_u1_u4_n118 ) , .ZN( u1_u1_u4_n131 ) , .A1( u1_u1_u4_n147 ) );
  NAND2_X1 u1_u1_u4_U22 (.A1( u1_u1_u4_n119 ) , .A2( u1_u1_u4_n120 ) , .ZN( u1_u1_u4_n130 ) );
  NAND2_X1 u1_u1_u4_U23 (.ZN( u1_u1_u4_n117 ) , .A2( u1_u1_u4_n118 ) , .A1( u1_u1_u4_n148 ) );
  NAND2_X1 u1_u1_u4_U24 (.ZN( u1_u1_u4_n129 ) , .A1( u1_u1_u4_n134 ) , .A2( u1_u1_u4_n148 ) );
  AND3_X1 u1_u1_u4_U25 (.A1( u1_u1_u4_n119 ) , .A2( u1_u1_u4_n143 ) , .A3( u1_u1_u4_n154 ) , .ZN( u1_u1_u4_n161 ) );
  AND2_X1 u1_u1_u4_U26 (.A1( u1_u1_u4_n145 ) , .A2( u1_u1_u4_n147 ) , .ZN( u1_u1_u4_n159 ) );
  OR3_X1 u1_u1_u4_U27 (.A3( u1_u1_u4_n114 ) , .A2( u1_u1_u4_n115 ) , .A1( u1_u1_u4_n116 ) , .ZN( u1_u1_u4_n136 ) );
  AOI21_X1 u1_u1_u4_U28 (.A( u1_u1_u4_n113 ) , .ZN( u1_u1_u4_n116 ) , .B2( u1_u1_u4_n173 ) , .B1( u1_u1_u4_n174 ) );
  AOI21_X1 u1_u1_u4_U29 (.ZN( u1_u1_u4_n115 ) , .B2( u1_u1_u4_n145 ) , .B1( u1_u1_u4_n146 ) , .A( u1_u1_u4_n156 ) );
  NOR2_X1 u1_u1_u4_U3 (.ZN( u1_u1_u4_n121 ) , .A1( u1_u1_u4_n181 ) , .A2( u1_u1_u4_n182 ) );
  OAI22_X1 u1_u1_u4_U30 (.ZN( u1_u1_u4_n114 ) , .A2( u1_u1_u4_n121 ) , .B1( u1_u1_u4_n160 ) , .B2( u1_u1_u4_n170 ) , .A1( u1_u1_u4_n171 ) );
  INV_X1 u1_u1_u4_U31 (.A( u1_u1_u4_n158 ) , .ZN( u1_u1_u4_n182 ) );
  INV_X1 u1_u1_u4_U32 (.ZN( u1_u1_u4_n181 ) , .A( u1_u1_u4_n96 ) );
  INV_X1 u1_u1_u4_U33 (.A( u1_u1_u4_n144 ) , .ZN( u1_u1_u4_n179 ) );
  INV_X1 u1_u1_u4_U34 (.A( u1_u1_u4_n157 ) , .ZN( u1_u1_u4_n178 ) );
  NAND2_X1 u1_u1_u4_U35 (.A2( u1_u1_u4_n154 ) , .A1( u1_u1_u4_n96 ) , .ZN( u1_u1_u4_n97 ) );
  INV_X1 u1_u1_u4_U36 (.ZN( u1_u1_u4_n186 ) , .A( u1_u1_u4_n95 ) );
  OAI221_X1 u1_u1_u4_U37 (.C1( u1_u1_u4_n134 ) , .B1( u1_u1_u4_n158 ) , .B2( u1_u1_u4_n171 ) , .C2( u1_u1_u4_n173 ) , .A( u1_u1_u4_n94 ) , .ZN( u1_u1_u4_n95 ) );
  AOI222_X1 u1_u1_u4_U38 (.B2( u1_u1_u4_n132 ) , .A1( u1_u1_u4_n138 ) , .C2( u1_u1_u4_n175 ) , .A2( u1_u1_u4_n179 ) , .C1( u1_u1_u4_n181 ) , .B1( u1_u1_u4_n185 ) , .ZN( u1_u1_u4_n94 ) );
  INV_X1 u1_u1_u4_U39 (.A( u1_u1_u4_n113 ) , .ZN( u1_u1_u4_n185 ) );
  INV_X1 u1_u1_u4_U4 (.A( u1_u1_u4_n117 ) , .ZN( u1_u1_u4_n184 ) );
  INV_X1 u1_u1_u4_U40 (.A( u1_u1_u4_n143 ) , .ZN( u1_u1_u4_n183 ) );
  NOR2_X1 u1_u1_u4_U41 (.ZN( u1_u1_u4_n138 ) , .A1( u1_u1_u4_n168 ) , .A2( u1_u1_u4_n169 ) );
  NOR2_X1 u1_u1_u4_U42 (.A1( u1_u1_u4_n150 ) , .A2( u1_u1_u4_n152 ) , .ZN( u1_u1_u4_n153 ) );
  NOR2_X1 u1_u1_u4_U43 (.A2( u1_u1_u4_n128 ) , .A1( u1_u1_u4_n138 ) , .ZN( u1_u1_u4_n156 ) );
  AOI22_X1 u1_u1_u4_U44 (.B2( u1_u1_u4_n122 ) , .A1( u1_u1_u4_n123 ) , .ZN( u1_u1_u4_n124 ) , .B1( u1_u1_u4_n128 ) , .A2( u1_u1_u4_n172 ) );
  NAND2_X1 u1_u1_u4_U45 (.A2( u1_u1_u4_n120 ) , .ZN( u1_u1_u4_n123 ) , .A1( u1_u1_u4_n161 ) );
  INV_X1 u1_u1_u4_U46 (.A( u1_u1_u4_n153 ) , .ZN( u1_u1_u4_n172 ) );
  AOI22_X1 u1_u1_u4_U47 (.B2( u1_u1_u4_n132 ) , .A2( u1_u1_u4_n133 ) , .ZN( u1_u1_u4_n140 ) , .A1( u1_u1_u4_n150 ) , .B1( u1_u1_u4_n179 ) );
  NAND2_X1 u1_u1_u4_U48 (.ZN( u1_u1_u4_n133 ) , .A2( u1_u1_u4_n146 ) , .A1( u1_u1_u4_n154 ) );
  NAND2_X1 u1_u1_u4_U49 (.A1( u1_u1_u4_n103 ) , .ZN( u1_u1_u4_n154 ) , .A2( u1_u1_u4_n98 ) );
  NOR4_X1 u1_u1_u4_U5 (.A4( u1_u1_u4_n106 ) , .A3( u1_u1_u4_n107 ) , .A2( u1_u1_u4_n108 ) , .A1( u1_u1_u4_n109 ) , .ZN( u1_u1_u4_n110 ) );
  NAND2_X1 u1_u1_u4_U50 (.A1( u1_u1_u4_n101 ) , .ZN( u1_u1_u4_n158 ) , .A2( u1_u1_u4_n99 ) );
  AOI21_X1 u1_u1_u4_U51 (.ZN( u1_u1_u4_n127 ) , .A( u1_u1_u4_n136 ) , .B2( u1_u1_u4_n150 ) , .B1( u1_u1_u4_n180 ) );
  INV_X1 u1_u1_u4_U52 (.A( u1_u1_u4_n160 ) , .ZN( u1_u1_u4_n180 ) );
  NAND2_X1 u1_u1_u4_U53 (.A2( u1_u1_u4_n104 ) , .A1( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n146 ) );
  NAND2_X1 u1_u1_u4_U54 (.A2( u1_u1_u4_n101 ) , .A1( u1_u1_u4_n102 ) , .ZN( u1_u1_u4_n160 ) );
  NAND2_X1 u1_u1_u4_U55 (.ZN( u1_u1_u4_n134 ) , .A1( u1_u1_u4_n98 ) , .A2( u1_u1_u4_n99 ) );
  NAND2_X1 u1_u1_u4_U56 (.A1( u1_u1_u4_n103 ) , .A2( u1_u1_u4_n104 ) , .ZN( u1_u1_u4_n143 ) );
  NAND2_X1 u1_u1_u4_U57 (.A2( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n145 ) , .A1( u1_u1_u4_n98 ) );
  NAND2_X1 u1_u1_u4_U58 (.A1( u1_u1_u4_n100 ) , .A2( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n120 ) );
  NAND2_X1 u1_u1_u4_U59 (.A1( u1_u1_u4_n102 ) , .A2( u1_u1_u4_n104 ) , .ZN( u1_u1_u4_n148 ) );
  AOI21_X1 u1_u1_u4_U6 (.ZN( u1_u1_u4_n106 ) , .B2( u1_u1_u4_n146 ) , .B1( u1_u1_u4_n158 ) , .A( u1_u1_u4_n170 ) );
  NAND2_X1 u1_u1_u4_U60 (.A2( u1_u1_u4_n100 ) , .A1( u1_u1_u4_n103 ) , .ZN( u1_u1_u4_n157 ) );
  INV_X1 u1_u1_u4_U61 (.A( u1_u1_u4_n150 ) , .ZN( u1_u1_u4_n173 ) );
  INV_X1 u1_u1_u4_U62 (.A( u1_u1_u4_n152 ) , .ZN( u1_u1_u4_n171 ) );
  NAND2_X1 u1_u1_u4_U63 (.A1( u1_u1_u4_n100 ) , .ZN( u1_u1_u4_n118 ) , .A2( u1_u1_u4_n99 ) );
  NAND2_X1 u1_u1_u4_U64 (.A2( u1_u1_u4_n100 ) , .A1( u1_u1_u4_n102 ) , .ZN( u1_u1_u4_n144 ) );
  NAND2_X1 u1_u1_u4_U65 (.A2( u1_u1_u4_n101 ) , .A1( u1_u1_u4_n105 ) , .ZN( u1_u1_u4_n96 ) );
  INV_X1 u1_u1_u4_U66 (.A( u1_u1_u4_n128 ) , .ZN( u1_u1_u4_n174 ) );
  NAND2_X1 u1_u1_u4_U67 (.A2( u1_u1_u4_n102 ) , .ZN( u1_u1_u4_n119 ) , .A1( u1_u1_u4_n98 ) );
  NAND2_X1 u1_u1_u4_U68 (.A2( u1_u1_u4_n101 ) , .A1( u1_u1_u4_n103 ) , .ZN( u1_u1_u4_n147 ) );
  NAND2_X1 u1_u1_u4_U69 (.A2( u1_u1_u4_n104 ) , .ZN( u1_u1_u4_n113 ) , .A1( u1_u1_u4_n99 ) );
  AOI21_X1 u1_u1_u4_U7 (.ZN( u1_u1_u4_n108 ) , .B2( u1_u1_u4_n134 ) , .B1( u1_u1_u4_n155 ) , .A( u1_u1_u4_n156 ) );
  NOR2_X1 u1_u1_u4_U70 (.A2( u1_u1_X_28 ) , .ZN( u1_u1_u4_n150 ) , .A1( u1_u1_u4_n168 ) );
  NOR2_X1 u1_u1_u4_U71 (.A2( u1_u1_X_29 ) , .ZN( u1_u1_u4_n152 ) , .A1( u1_u1_u4_n169 ) );
  NOR2_X1 u1_u1_u4_U72 (.A2( u1_u1_X_30 ) , .ZN( u1_u1_u4_n105 ) , .A1( u1_u1_u4_n176 ) );
  NOR2_X1 u1_u1_u4_U73 (.A2( u1_u1_X_26 ) , .ZN( u1_u1_u4_n100 ) , .A1( u1_u1_u4_n177 ) );
  NOR2_X1 u1_u1_u4_U74 (.A2( u1_u1_X_28 ) , .A1( u1_u1_X_29 ) , .ZN( u1_u1_u4_n128 ) );
  NOR2_X1 u1_u1_u4_U75 (.A2( u1_u1_X_27 ) , .A1( u1_u1_X_30 ) , .ZN( u1_u1_u4_n102 ) );
  NOR2_X1 u1_u1_u4_U76 (.A2( u1_u1_X_25 ) , .A1( u1_u1_X_26 ) , .ZN( u1_u1_u4_n98 ) );
  AND2_X1 u1_u1_u4_U77 (.A2( u1_u1_X_25 ) , .A1( u1_u1_X_26 ) , .ZN( u1_u1_u4_n104 ) );
  AND2_X1 u1_u1_u4_U78 (.A1( u1_u1_X_30 ) , .A2( u1_u1_u4_n176 ) , .ZN( u1_u1_u4_n99 ) );
  AND2_X1 u1_u1_u4_U79 (.A1( u1_u1_X_26 ) , .ZN( u1_u1_u4_n101 ) , .A2( u1_u1_u4_n177 ) );
  AOI21_X1 u1_u1_u4_U8 (.ZN( u1_u1_u4_n109 ) , .A( u1_u1_u4_n153 ) , .B1( u1_u1_u4_n159 ) , .B2( u1_u1_u4_n184 ) );
  AND2_X1 u1_u1_u4_U80 (.A1( u1_u1_X_27 ) , .A2( u1_u1_X_30 ) , .ZN( u1_u1_u4_n103 ) );
  INV_X1 u1_u1_u4_U81 (.A( u1_u1_X_28 ) , .ZN( u1_u1_u4_n169 ) );
  INV_X1 u1_u1_u4_U82 (.A( u1_u1_X_29 ) , .ZN( u1_u1_u4_n168 ) );
  INV_X1 u1_u1_u4_U83 (.A( u1_u1_X_25 ) , .ZN( u1_u1_u4_n177 ) );
  INV_X1 u1_u1_u4_U84 (.A( u1_u1_X_27 ) , .ZN( u1_u1_u4_n176 ) );
  NAND4_X1 u1_u1_u4_U85 (.ZN( u1_out1_25 ) , .A4( u1_u1_u4_n139 ) , .A3( u1_u1_u4_n140 ) , .A2( u1_u1_u4_n141 ) , .A1( u1_u1_u4_n142 ) );
  OAI21_X1 u1_u1_u4_U86 (.A( u1_u1_u4_n128 ) , .B2( u1_u1_u4_n129 ) , .B1( u1_u1_u4_n130 ) , .ZN( u1_u1_u4_n142 ) );
  OAI21_X1 u1_u1_u4_U87 (.B2( u1_u1_u4_n131 ) , .ZN( u1_u1_u4_n141 ) , .A( u1_u1_u4_n175 ) , .B1( u1_u1_u4_n183 ) );
  NAND4_X1 u1_u1_u4_U88 (.ZN( u1_out1_14 ) , .A4( u1_u1_u4_n124 ) , .A3( u1_u1_u4_n125 ) , .A2( u1_u1_u4_n126 ) , .A1( u1_u1_u4_n127 ) );
  AOI22_X1 u1_u1_u4_U89 (.B2( u1_u1_u4_n117 ) , .ZN( u1_u1_u4_n126 ) , .A1( u1_u1_u4_n129 ) , .B1( u1_u1_u4_n152 ) , .A2( u1_u1_u4_n175 ) );
  AOI211_X1 u1_u1_u4_U9 (.B( u1_u1_u4_n136 ) , .A( u1_u1_u4_n137 ) , .C2( u1_u1_u4_n138 ) , .ZN( u1_u1_u4_n139 ) , .C1( u1_u1_u4_n182 ) );
  AOI22_X1 u1_u1_u4_U90 (.ZN( u1_u1_u4_n125 ) , .B2( u1_u1_u4_n131 ) , .A2( u1_u1_u4_n132 ) , .B1( u1_u1_u4_n138 ) , .A1( u1_u1_u4_n178 ) );
  NAND4_X1 u1_u1_u4_U91 (.ZN( u1_out1_8 ) , .A4( u1_u1_u4_n110 ) , .A3( u1_u1_u4_n111 ) , .A2( u1_u1_u4_n112 ) , .A1( u1_u1_u4_n186 ) );
  NAND2_X1 u1_u1_u4_U92 (.ZN( u1_u1_u4_n112 ) , .A2( u1_u1_u4_n130 ) , .A1( u1_u1_u4_n150 ) );
  AOI22_X1 u1_u1_u4_U93 (.ZN( u1_u1_u4_n111 ) , .B2( u1_u1_u4_n132 ) , .A1( u1_u1_u4_n152 ) , .B1( u1_u1_u4_n178 ) , .A2( u1_u1_u4_n97 ) );
  AOI22_X1 u1_u1_u4_U94 (.B2( u1_u1_u4_n149 ) , .B1( u1_u1_u4_n150 ) , .A2( u1_u1_u4_n151 ) , .A1( u1_u1_u4_n152 ) , .ZN( u1_u1_u4_n167 ) );
  NOR4_X1 u1_u1_u4_U95 (.A4( u1_u1_u4_n162 ) , .A3( u1_u1_u4_n163 ) , .A2( u1_u1_u4_n164 ) , .A1( u1_u1_u4_n165 ) , .ZN( u1_u1_u4_n166 ) );
  NAND3_X1 u1_u1_u4_U96 (.ZN( u1_out1_3 ) , .A3( u1_u1_u4_n166 ) , .A1( u1_u1_u4_n167 ) , .A2( u1_u1_u4_n186 ) );
  NAND3_X1 u1_u1_u4_U97 (.A3( u1_u1_u4_n146 ) , .A2( u1_u1_u4_n147 ) , .A1( u1_u1_u4_n148 ) , .ZN( u1_u1_u4_n149 ) );
  NAND3_X1 u1_u1_u4_U98 (.A3( u1_u1_u4_n143 ) , .A2( u1_u1_u4_n144 ) , .A1( u1_u1_u4_n145 ) , .ZN( u1_u1_u4_n151 ) );
  NAND3_X1 u1_u1_u4_U99 (.A3( u1_u1_u4_n121 ) , .ZN( u1_u1_u4_n122 ) , .A2( u1_u1_u4_n144 ) , .A1( u1_u1_u4_n154 ) );
  AOI22_X1 u1_u1_u6_U10 (.A2( u1_u1_u6_n151 ) , .B2( u1_u1_u6_n161 ) , .A1( u1_u1_u6_n167 ) , .B1( u1_u1_u6_n170 ) , .ZN( u1_u1_u6_n89 ) );
  AOI21_X1 u1_u1_u6_U11 (.B1( u1_u1_u6_n107 ) , .B2( u1_u1_u6_n132 ) , .A( u1_u1_u6_n158 ) , .ZN( u1_u1_u6_n88 ) );
  AOI21_X1 u1_u1_u6_U12 (.B2( u1_u1_u6_n147 ) , .B1( u1_u1_u6_n148 ) , .ZN( u1_u1_u6_n149 ) , .A( u1_u1_u6_n158 ) );
  AOI21_X1 u1_u1_u6_U13 (.ZN( u1_u1_u6_n106 ) , .A( u1_u1_u6_n142 ) , .B2( u1_u1_u6_n159 ) , .B1( u1_u1_u6_n164 ) );
  INV_X1 u1_u1_u6_U14 (.A( u1_u1_u6_n155 ) , .ZN( u1_u1_u6_n161 ) );
  INV_X1 u1_u1_u6_U15 (.A( u1_u1_u6_n128 ) , .ZN( u1_u1_u6_n164 ) );
  NAND2_X1 u1_u1_u6_U16 (.ZN( u1_u1_u6_n110 ) , .A1( u1_u1_u6_n122 ) , .A2( u1_u1_u6_n129 ) );
  NAND2_X1 u1_u1_u6_U17 (.ZN( u1_u1_u6_n124 ) , .A2( u1_u1_u6_n146 ) , .A1( u1_u1_u6_n148 ) );
  INV_X1 u1_u1_u6_U18 (.A( u1_u1_u6_n132 ) , .ZN( u1_u1_u6_n171 ) );
  AND2_X1 u1_u1_u6_U19 (.A1( u1_u1_u6_n100 ) , .ZN( u1_u1_u6_n130 ) , .A2( u1_u1_u6_n147 ) );
  INV_X1 u1_u1_u6_U20 (.A( u1_u1_u6_n127 ) , .ZN( u1_u1_u6_n173 ) );
  INV_X1 u1_u1_u6_U21 (.A( u1_u1_u6_n121 ) , .ZN( u1_u1_u6_n167 ) );
  INV_X1 u1_u1_u6_U22 (.A( u1_u1_u6_n100 ) , .ZN( u1_u1_u6_n169 ) );
  INV_X1 u1_u1_u6_U23 (.A( u1_u1_u6_n123 ) , .ZN( u1_u1_u6_n170 ) );
  INV_X1 u1_u1_u6_U24 (.A( u1_u1_u6_n113 ) , .ZN( u1_u1_u6_n168 ) );
  AND2_X1 u1_u1_u6_U25 (.A1( u1_u1_u6_n107 ) , .A2( u1_u1_u6_n119 ) , .ZN( u1_u1_u6_n133 ) );
  AND2_X1 u1_u1_u6_U26 (.A2( u1_u1_u6_n121 ) , .A1( u1_u1_u6_n122 ) , .ZN( u1_u1_u6_n131 ) );
  AND3_X1 u1_u1_u6_U27 (.ZN( u1_u1_u6_n120 ) , .A2( u1_u1_u6_n127 ) , .A1( u1_u1_u6_n132 ) , .A3( u1_u1_u6_n145 ) );
  INV_X1 u1_u1_u6_U28 (.A( u1_u1_u6_n146 ) , .ZN( u1_u1_u6_n163 ) );
  AOI222_X1 u1_u1_u6_U29 (.ZN( u1_u1_u6_n114 ) , .A1( u1_u1_u6_n118 ) , .A2( u1_u1_u6_n126 ) , .B2( u1_u1_u6_n151 ) , .C2( u1_u1_u6_n159 ) , .C1( u1_u1_u6_n168 ) , .B1( u1_u1_u6_n169 ) );
  INV_X1 u1_u1_u6_U3 (.A( u1_u1_u6_n110 ) , .ZN( u1_u1_u6_n166 ) );
  NOR2_X1 u1_u1_u6_U30 (.A1( u1_u1_u6_n162 ) , .A2( u1_u1_u6_n165 ) , .ZN( u1_u1_u6_n98 ) );
  AOI211_X1 u1_u1_u6_U31 (.B( u1_u1_u6_n134 ) , .A( u1_u1_u6_n135 ) , .C1( u1_u1_u6_n136 ) , .ZN( u1_u1_u6_n137 ) , .C2( u1_u1_u6_n151 ) );
  AOI21_X1 u1_u1_u6_U32 (.B1( u1_u1_u6_n131 ) , .ZN( u1_u1_u6_n135 ) , .A( u1_u1_u6_n144 ) , .B2( u1_u1_u6_n146 ) );
  NAND4_X1 u1_u1_u6_U33 (.A4( u1_u1_u6_n127 ) , .A3( u1_u1_u6_n128 ) , .A2( u1_u1_u6_n129 ) , .A1( u1_u1_u6_n130 ) , .ZN( u1_u1_u6_n136 ) );
  AOI21_X1 u1_u1_u6_U34 (.B2( u1_u1_u6_n132 ) , .B1( u1_u1_u6_n133 ) , .ZN( u1_u1_u6_n134 ) , .A( u1_u1_u6_n158 ) );
  NAND2_X1 u1_u1_u6_U35 (.A1( u1_u1_u6_n144 ) , .ZN( u1_u1_u6_n151 ) , .A2( u1_u1_u6_n158 ) );
  NAND2_X1 u1_u1_u6_U36 (.ZN( u1_u1_u6_n132 ) , .A1( u1_u1_u6_n91 ) , .A2( u1_u1_u6_n97 ) );
  AOI22_X1 u1_u1_u6_U37 (.B2( u1_u1_u6_n110 ) , .B1( u1_u1_u6_n111 ) , .A1( u1_u1_u6_n112 ) , .ZN( u1_u1_u6_n115 ) , .A2( u1_u1_u6_n161 ) );
  NAND4_X1 u1_u1_u6_U38 (.A3( u1_u1_u6_n109 ) , .ZN( u1_u1_u6_n112 ) , .A4( u1_u1_u6_n132 ) , .A2( u1_u1_u6_n147 ) , .A1( u1_u1_u6_n166 ) );
  NOR2_X1 u1_u1_u6_U39 (.ZN( u1_u1_u6_n109 ) , .A1( u1_u1_u6_n170 ) , .A2( u1_u1_u6_n173 ) );
  INV_X1 u1_u1_u6_U4 (.A( u1_u1_u6_n142 ) , .ZN( u1_u1_u6_n174 ) );
  NOR2_X1 u1_u1_u6_U40 (.A2( u1_u1_u6_n126 ) , .ZN( u1_u1_u6_n155 ) , .A1( u1_u1_u6_n160 ) );
  NAND2_X1 u1_u1_u6_U41 (.ZN( u1_u1_u6_n146 ) , .A2( u1_u1_u6_n94 ) , .A1( u1_u1_u6_n99 ) );
  AOI21_X1 u1_u1_u6_U42 (.A( u1_u1_u6_n144 ) , .B2( u1_u1_u6_n145 ) , .B1( u1_u1_u6_n146 ) , .ZN( u1_u1_u6_n150 ) );
  INV_X1 u1_u1_u6_U43 (.A( u1_u1_u6_n111 ) , .ZN( u1_u1_u6_n158 ) );
  NAND2_X1 u1_u1_u6_U44 (.ZN( u1_u1_u6_n127 ) , .A1( u1_u1_u6_n91 ) , .A2( u1_u1_u6_n92 ) );
  NAND2_X1 u1_u1_u6_U45 (.ZN( u1_u1_u6_n129 ) , .A2( u1_u1_u6_n95 ) , .A1( u1_u1_u6_n96 ) );
  INV_X1 u1_u1_u6_U46 (.A( u1_u1_u6_n144 ) , .ZN( u1_u1_u6_n159 ) );
  NAND2_X1 u1_u1_u6_U47 (.ZN( u1_u1_u6_n145 ) , .A2( u1_u1_u6_n97 ) , .A1( u1_u1_u6_n98 ) );
  NAND2_X1 u1_u1_u6_U48 (.ZN( u1_u1_u6_n148 ) , .A2( u1_u1_u6_n92 ) , .A1( u1_u1_u6_n94 ) );
  NAND2_X1 u1_u1_u6_U49 (.ZN( u1_u1_u6_n108 ) , .A2( u1_u1_u6_n139 ) , .A1( u1_u1_u6_n144 ) );
  NAND2_X1 u1_u1_u6_U5 (.A2( u1_u1_u6_n143 ) , .ZN( u1_u1_u6_n152 ) , .A1( u1_u1_u6_n166 ) );
  NAND2_X1 u1_u1_u6_U50 (.ZN( u1_u1_u6_n121 ) , .A2( u1_u1_u6_n95 ) , .A1( u1_u1_u6_n97 ) );
  NAND2_X1 u1_u1_u6_U51 (.ZN( u1_u1_u6_n107 ) , .A2( u1_u1_u6_n92 ) , .A1( u1_u1_u6_n95 ) );
  AND2_X1 u1_u1_u6_U52 (.ZN( u1_u1_u6_n118 ) , .A2( u1_u1_u6_n91 ) , .A1( u1_u1_u6_n99 ) );
  NAND2_X1 u1_u1_u6_U53 (.ZN( u1_u1_u6_n147 ) , .A2( u1_u1_u6_n98 ) , .A1( u1_u1_u6_n99 ) );
  NAND2_X1 u1_u1_u6_U54 (.ZN( u1_u1_u6_n128 ) , .A1( u1_u1_u6_n94 ) , .A2( u1_u1_u6_n96 ) );
  NAND2_X1 u1_u1_u6_U55 (.ZN( u1_u1_u6_n119 ) , .A2( u1_u1_u6_n95 ) , .A1( u1_u1_u6_n99 ) );
  NAND2_X1 u1_u1_u6_U56 (.ZN( u1_u1_u6_n123 ) , .A2( u1_u1_u6_n91 ) , .A1( u1_u1_u6_n96 ) );
  NAND2_X1 u1_u1_u6_U57 (.ZN( u1_u1_u6_n100 ) , .A2( u1_u1_u6_n92 ) , .A1( u1_u1_u6_n98 ) );
  NAND2_X1 u1_u1_u6_U58 (.ZN( u1_u1_u6_n122 ) , .A1( u1_u1_u6_n94 ) , .A2( u1_u1_u6_n97 ) );
  INV_X1 u1_u1_u6_U59 (.A( u1_u1_u6_n139 ) , .ZN( u1_u1_u6_n160 ) );
  AOI22_X1 u1_u1_u6_U6 (.B2( u1_u1_u6_n101 ) , .A1( u1_u1_u6_n102 ) , .ZN( u1_u1_u6_n103 ) , .B1( u1_u1_u6_n160 ) , .A2( u1_u1_u6_n161 ) );
  NAND2_X1 u1_u1_u6_U60 (.ZN( u1_u1_u6_n113 ) , .A1( u1_u1_u6_n96 ) , .A2( u1_u1_u6_n98 ) );
  NOR2_X1 u1_u1_u6_U61 (.A2( u1_u1_X_40 ) , .A1( u1_u1_X_41 ) , .ZN( u1_u1_u6_n126 ) );
  NOR2_X1 u1_u1_u6_U62 (.A2( u1_u1_X_39 ) , .A1( u1_u1_X_42 ) , .ZN( u1_u1_u6_n92 ) );
  NOR2_X1 u1_u1_u6_U63 (.A2( u1_u1_X_39 ) , .A1( u1_u1_u6_n156 ) , .ZN( u1_u1_u6_n97 ) );
  NOR2_X1 u1_u1_u6_U64 (.A2( u1_u1_X_38 ) , .A1( u1_u1_u6_n165 ) , .ZN( u1_u1_u6_n95 ) );
  NOR2_X1 u1_u1_u6_U65 (.A2( u1_u1_X_41 ) , .ZN( u1_u1_u6_n111 ) , .A1( u1_u1_u6_n157 ) );
  NOR2_X1 u1_u1_u6_U66 (.A2( u1_u1_X_37 ) , .A1( u1_u1_u6_n162 ) , .ZN( u1_u1_u6_n94 ) );
  NOR2_X1 u1_u1_u6_U67 (.A2( u1_u1_X_37 ) , .A1( u1_u1_X_38 ) , .ZN( u1_u1_u6_n91 ) );
  NAND2_X1 u1_u1_u6_U68 (.A1( u1_u1_X_41 ) , .ZN( u1_u1_u6_n144 ) , .A2( u1_u1_u6_n157 ) );
  NAND2_X1 u1_u1_u6_U69 (.A2( u1_u1_X_40 ) , .A1( u1_u1_X_41 ) , .ZN( u1_u1_u6_n139 ) );
  NOR2_X1 u1_u1_u6_U7 (.A1( u1_u1_u6_n118 ) , .ZN( u1_u1_u6_n143 ) , .A2( u1_u1_u6_n168 ) );
  AND2_X1 u1_u1_u6_U70 (.A1( u1_u1_X_39 ) , .A2( u1_u1_u6_n156 ) , .ZN( u1_u1_u6_n96 ) );
  AND2_X1 u1_u1_u6_U71 (.A1( u1_u1_X_39 ) , .A2( u1_u1_X_42 ) , .ZN( u1_u1_u6_n99 ) );
  INV_X1 u1_u1_u6_U72 (.A( u1_u1_X_40 ) , .ZN( u1_u1_u6_n157 ) );
  INV_X1 u1_u1_u6_U73 (.A( u1_u1_X_37 ) , .ZN( u1_u1_u6_n165 ) );
  INV_X1 u1_u1_u6_U74 (.A( u1_u1_X_38 ) , .ZN( u1_u1_u6_n162 ) );
  INV_X1 u1_u1_u6_U75 (.A( u1_u1_X_42 ) , .ZN( u1_u1_u6_n156 ) );
  NAND4_X1 u1_u1_u6_U76 (.ZN( u1_out1_32 ) , .A4( u1_u1_u6_n103 ) , .A3( u1_u1_u6_n104 ) , .A2( u1_u1_u6_n105 ) , .A1( u1_u1_u6_n106 ) );
  AOI22_X1 u1_u1_u6_U77 (.ZN( u1_u1_u6_n105 ) , .A2( u1_u1_u6_n108 ) , .A1( u1_u1_u6_n118 ) , .B2( u1_u1_u6_n126 ) , .B1( u1_u1_u6_n171 ) );
  AOI22_X1 u1_u1_u6_U78 (.ZN( u1_u1_u6_n104 ) , .A1( u1_u1_u6_n111 ) , .B1( u1_u1_u6_n124 ) , .B2( u1_u1_u6_n151 ) , .A2( u1_u1_u6_n93 ) );
  NAND4_X1 u1_u1_u6_U79 (.ZN( u1_out1_12 ) , .A4( u1_u1_u6_n114 ) , .A3( u1_u1_u6_n115 ) , .A2( u1_u1_u6_n116 ) , .A1( u1_u1_u6_n117 ) );
  OAI21_X1 u1_u1_u6_U8 (.A( u1_u1_u6_n159 ) , .B1( u1_u1_u6_n169 ) , .B2( u1_u1_u6_n173 ) , .ZN( u1_u1_u6_n90 ) );
  OAI22_X1 u1_u1_u6_U80 (.B2( u1_u1_u6_n111 ) , .ZN( u1_u1_u6_n116 ) , .B1( u1_u1_u6_n126 ) , .A2( u1_u1_u6_n164 ) , .A1( u1_u1_u6_n167 ) );
  OAI21_X1 u1_u1_u6_U81 (.A( u1_u1_u6_n108 ) , .ZN( u1_u1_u6_n117 ) , .B2( u1_u1_u6_n141 ) , .B1( u1_u1_u6_n163 ) );
  OAI211_X1 u1_u1_u6_U82 (.ZN( u1_out1_7 ) , .B( u1_u1_u6_n153 ) , .C2( u1_u1_u6_n154 ) , .C1( u1_u1_u6_n155 ) , .A( u1_u1_u6_n174 ) );
  NOR3_X1 u1_u1_u6_U83 (.A1( u1_u1_u6_n141 ) , .ZN( u1_u1_u6_n154 ) , .A3( u1_u1_u6_n164 ) , .A2( u1_u1_u6_n171 ) );
  AOI211_X1 u1_u1_u6_U84 (.B( u1_u1_u6_n149 ) , .A( u1_u1_u6_n150 ) , .C2( u1_u1_u6_n151 ) , .C1( u1_u1_u6_n152 ) , .ZN( u1_u1_u6_n153 ) );
  OAI211_X1 u1_u1_u6_U85 (.ZN( u1_out1_22 ) , .B( u1_u1_u6_n137 ) , .A( u1_u1_u6_n138 ) , .C2( u1_u1_u6_n139 ) , .C1( u1_u1_u6_n140 ) );
  AND4_X1 u1_u1_u6_U86 (.A3( u1_u1_u6_n119 ) , .A1( u1_u1_u6_n120 ) , .A4( u1_u1_u6_n129 ) , .ZN( u1_u1_u6_n140 ) , .A2( u1_u1_u6_n143 ) );
  AOI22_X1 u1_u1_u6_U87 (.B1( u1_u1_u6_n124 ) , .A2( u1_u1_u6_n125 ) , .A1( u1_u1_u6_n126 ) , .ZN( u1_u1_u6_n138 ) , .B2( u1_u1_u6_n161 ) );
  NAND3_X1 u1_u1_u6_U88 (.A2( u1_u1_u6_n123 ) , .ZN( u1_u1_u6_n125 ) , .A1( u1_u1_u6_n130 ) , .A3( u1_u1_u6_n131 ) );
  NAND3_X1 u1_u1_u6_U89 (.A3( u1_u1_u6_n133 ) , .ZN( u1_u1_u6_n141 ) , .A1( u1_u1_u6_n145 ) , .A2( u1_u1_u6_n148 ) );
  INV_X1 u1_u1_u6_U9 (.ZN( u1_u1_u6_n172 ) , .A( u1_u1_u6_n88 ) );
  NAND3_X1 u1_u1_u6_U90 (.ZN( u1_u1_u6_n101 ) , .A3( u1_u1_u6_n107 ) , .A2( u1_u1_u6_n121 ) , .A1( u1_u1_u6_n127 ) );
  NAND3_X1 u1_u1_u6_U91 (.ZN( u1_u1_u6_n102 ) , .A3( u1_u1_u6_n130 ) , .A2( u1_u1_u6_n145 ) , .A1( u1_u1_u6_n166 ) );
  NAND3_X1 u1_u1_u6_U92 (.A3( u1_u1_u6_n113 ) , .A1( u1_u1_u6_n119 ) , .A2( u1_u1_u6_n123 ) , .ZN( u1_u1_u6_n93 ) );
  NAND3_X1 u1_u1_u6_U93 (.ZN( u1_u1_u6_n142 ) , .A2( u1_u1_u6_n172 ) , .A3( u1_u1_u6_n89 ) , .A1( u1_u1_u6_n90 ) );
  XOR2_X1 u1_u2_U1 (.B( u1_K3_9 ) , .A( u1_R1_6 ) , .Z( u1_u2_X_9 ) );
  XOR2_X1 u1_u2_U16 (.B( u1_K3_3 ) , .A( u1_R1_2 ) , .Z( u1_u2_X_3 ) );
  XOR2_X1 u1_u2_U2 (.B( u1_K3_8 ) , .A( u1_R1_5 ) , .Z( u1_u2_X_8 ) );
  XOR2_X1 u1_u2_U27 (.B( u1_K3_2 ) , .A( u1_R1_1 ) , .Z( u1_u2_X_2 ) );
  XOR2_X1 u1_u2_U3 (.B( u1_K3_7 ) , .A( u1_R1_4 ) , .Z( u1_u2_X_7 ) );
  XOR2_X1 u1_u2_U33 (.B( u1_K3_24 ) , .A( u1_R1_17 ) , .Z( u1_u2_X_24 ) );
  XOR2_X1 u1_u2_U34 (.B( u1_K3_23 ) , .A( u1_R1_16 ) , .Z( u1_u2_X_23 ) );
  XOR2_X1 u1_u2_U35 (.B( u1_K3_22 ) , .A( u1_R1_15 ) , .Z( u1_u2_X_22 ) );
  XOR2_X1 u1_u2_U36 (.B( u1_K3_21 ) , .A( u1_R1_14 ) , .Z( u1_u2_X_21 ) );
  XOR2_X1 u1_u2_U37 (.B( u1_K3_20 ) , .A( u1_R1_13 ) , .Z( u1_u2_X_20 ) );
  XOR2_X1 u1_u2_U38 (.B( u1_K3_1 ) , .A( u1_R1_32 ) , .Z( u1_u2_X_1 ) );
  XOR2_X1 u1_u2_U39 (.B( u1_K3_19 ) , .A( u1_R1_12 ) , .Z( u1_u2_X_19 ) );
  XOR2_X1 u1_u2_U4 (.B( u1_K3_6 ) , .A( u1_R1_5 ) , .Z( u1_u2_X_6 ) );
  XOR2_X1 u1_u2_U40 (.B( u1_K3_18 ) , .A( u1_R1_13 ) , .Z( u1_u2_X_18 ) );
  XOR2_X1 u1_u2_U41 (.B( u1_K3_17 ) , .A( u1_R1_12 ) , .Z( u1_u2_X_17 ) );
  XOR2_X1 u1_u2_U42 (.B( u1_K3_16 ) , .A( u1_R1_11 ) , .Z( u1_u2_X_16 ) );
  XOR2_X1 u1_u2_U43 (.B( u1_K3_15 ) , .A( u1_R1_10 ) , .Z( u1_u2_X_15 ) );
  XOR2_X1 u1_u2_U44 (.B( u1_K3_14 ) , .A( u1_R1_9 ) , .Z( u1_u2_X_14 ) );
  XOR2_X1 u1_u2_U45 (.B( u1_K3_13 ) , .A( u1_R1_8 ) , .Z( u1_u2_X_13 ) );
  XOR2_X1 u1_u2_U46 (.B( u1_K3_12 ) , .A( u1_R1_9 ) , .Z( u1_u2_X_12 ) );
  XOR2_X1 u1_u2_U47 (.B( u1_K3_11 ) , .A( u1_R1_8 ) , .Z( u1_u2_X_11 ) );
  XOR2_X1 u1_u2_U48 (.B( u1_K3_10 ) , .A( u1_R1_7 ) , .Z( u1_u2_X_10 ) );
  XOR2_X1 u1_u2_U5 (.B( u1_K3_5 ) , .A( u1_R1_4 ) , .Z( u1_u2_X_5 ) );
  XOR2_X1 u1_u2_U6 (.B( u1_K3_4 ) , .A( u1_R1_3 ) , .Z( u1_u2_X_4 ) );
  AND3_X1 u1_u2_u0_U10 (.A2( u1_u2_u0_n112 ) , .ZN( u1_u2_u0_n127 ) , .A3( u1_u2_u0_n130 ) , .A1( u1_u2_u0_n148 ) );
  NAND2_X1 u1_u2_u0_U11 (.ZN( u1_u2_u0_n113 ) , .A1( u1_u2_u0_n139 ) , .A2( u1_u2_u0_n149 ) );
  AND2_X1 u1_u2_u0_U12 (.ZN( u1_u2_u0_n107 ) , .A1( u1_u2_u0_n130 ) , .A2( u1_u2_u0_n140 ) );
  AND2_X1 u1_u2_u0_U13 (.A2( u1_u2_u0_n129 ) , .A1( u1_u2_u0_n130 ) , .ZN( u1_u2_u0_n151 ) );
  AND2_X1 u1_u2_u0_U14 (.A1( u1_u2_u0_n108 ) , .A2( u1_u2_u0_n125 ) , .ZN( u1_u2_u0_n145 ) );
  INV_X1 u1_u2_u0_U15 (.A( u1_u2_u0_n143 ) , .ZN( u1_u2_u0_n173 ) );
  NOR2_X1 u1_u2_u0_U16 (.A2( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n147 ) , .A1( u1_u2_u0_n160 ) );
  INV_X1 u1_u2_u0_U17 (.ZN( u1_u2_u0_n172 ) , .A( u1_u2_u0_n88 ) );
  OAI222_X1 u1_u2_u0_U18 (.C1( u1_u2_u0_n108 ) , .A1( u1_u2_u0_n125 ) , .B2( u1_u2_u0_n128 ) , .B1( u1_u2_u0_n144 ) , .A2( u1_u2_u0_n158 ) , .C2( u1_u2_u0_n161 ) , .ZN( u1_u2_u0_n88 ) );
  NOR2_X1 u1_u2_u0_U19 (.A1( u1_u2_u0_n163 ) , .A2( u1_u2_u0_n164 ) , .ZN( u1_u2_u0_n95 ) );
  AOI21_X1 u1_u2_u0_U20 (.B1( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n132 ) , .A( u1_u2_u0_n165 ) , .B2( u1_u2_u0_n93 ) );
  INV_X1 u1_u2_u0_U21 (.A( u1_u2_u0_n142 ) , .ZN( u1_u2_u0_n165 ) );
  OAI221_X1 u1_u2_u0_U22 (.C1( u1_u2_u0_n121 ) , .ZN( u1_u2_u0_n122 ) , .B2( u1_u2_u0_n127 ) , .A( u1_u2_u0_n143 ) , .B1( u1_u2_u0_n144 ) , .C2( u1_u2_u0_n147 ) );
  OAI22_X1 u1_u2_u0_U23 (.B1( u1_u2_u0_n125 ) , .ZN( u1_u2_u0_n126 ) , .A1( u1_u2_u0_n138 ) , .A2( u1_u2_u0_n146 ) , .B2( u1_u2_u0_n147 ) );
  OAI22_X1 u1_u2_u0_U24 (.B1( u1_u2_u0_n131 ) , .A1( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n147 ) , .A2( u1_u2_u0_n90 ) , .ZN( u1_u2_u0_n91 ) );
  AND3_X1 u1_u2_u0_U25 (.A3( u1_u2_u0_n121 ) , .A2( u1_u2_u0_n125 ) , .A1( u1_u2_u0_n148 ) , .ZN( u1_u2_u0_n90 ) );
  INV_X1 u1_u2_u0_U26 (.A( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n161 ) );
  NOR2_X1 u1_u2_u0_U27 (.A1( u1_u2_u0_n120 ) , .ZN( u1_u2_u0_n143 ) , .A2( u1_u2_u0_n167 ) );
  OAI221_X1 u1_u2_u0_U28 (.C1( u1_u2_u0_n112 ) , .ZN( u1_u2_u0_n120 ) , .B1( u1_u2_u0_n138 ) , .B2( u1_u2_u0_n141 ) , .C2( u1_u2_u0_n147 ) , .A( u1_u2_u0_n172 ) );
  AOI211_X1 u1_u2_u0_U29 (.B( u1_u2_u0_n115 ) , .A( u1_u2_u0_n116 ) , .C2( u1_u2_u0_n117 ) , .C1( u1_u2_u0_n118 ) , .ZN( u1_u2_u0_n119 ) );
  INV_X1 u1_u2_u0_U3 (.A( u1_u2_u0_n113 ) , .ZN( u1_u2_u0_n166 ) );
  AOI22_X1 u1_u2_u0_U30 (.B2( u1_u2_u0_n109 ) , .A2( u1_u2_u0_n110 ) , .ZN( u1_u2_u0_n111 ) , .B1( u1_u2_u0_n118 ) , .A1( u1_u2_u0_n160 ) );
  INV_X1 u1_u2_u0_U31 (.A( u1_u2_u0_n118 ) , .ZN( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U32 (.ZN( u1_u2_u0_n104 ) , .B1( u1_u2_u0_n107 ) , .B2( u1_u2_u0_n141 ) , .A( u1_u2_u0_n144 ) );
  AOI21_X1 u1_u2_u0_U33 (.B1( u1_u2_u0_n127 ) , .B2( u1_u2_u0_n129 ) , .A( u1_u2_u0_n138 ) , .ZN( u1_u2_u0_n96 ) );
  AOI21_X1 u1_u2_u0_U34 (.ZN( u1_u2_u0_n116 ) , .B2( u1_u2_u0_n142 ) , .A( u1_u2_u0_n144 ) , .B1( u1_u2_u0_n166 ) );
  NAND2_X1 u1_u2_u0_U35 (.A1( u1_u2_u0_n100 ) , .A2( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n125 ) );
  NAND2_X1 u1_u2_u0_U36 (.A1( u1_u2_u0_n101 ) , .A2( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n150 ) );
  INV_X1 u1_u2_u0_U37 (.A( u1_u2_u0_n138 ) , .ZN( u1_u2_u0_n160 ) );
  NAND2_X1 u1_u2_u0_U38 (.A1( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n128 ) , .A2( u1_u2_u0_n95 ) );
  NAND2_X1 u1_u2_u0_U39 (.A1( u1_u2_u0_n100 ) , .ZN( u1_u2_u0_n129 ) , .A2( u1_u2_u0_n95 ) );
  AOI21_X1 u1_u2_u0_U4 (.B1( u1_u2_u0_n114 ) , .ZN( u1_u2_u0_n115 ) , .B2( u1_u2_u0_n129 ) , .A( u1_u2_u0_n161 ) );
  NAND2_X1 u1_u2_u0_U40 (.A2( u1_u2_u0_n100 ) , .ZN( u1_u2_u0_n131 ) , .A1( u1_u2_u0_n92 ) );
  NAND2_X1 u1_u2_u0_U41 (.A2( u1_u2_u0_n100 ) , .A1( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n139 ) );
  NAND2_X1 u1_u2_u0_U42 (.ZN( u1_u2_u0_n148 ) , .A1( u1_u2_u0_n93 ) , .A2( u1_u2_u0_n95 ) );
  NAND2_X1 u1_u2_u0_U43 (.A2( u1_u2_u0_n102 ) , .A1( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n149 ) );
  NAND2_X1 u1_u2_u0_U44 (.A2( u1_u2_u0_n102 ) , .ZN( u1_u2_u0_n114 ) , .A1( u1_u2_u0_n92 ) );
  NAND2_X1 u1_u2_u0_U45 (.A2( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n121 ) , .A1( u1_u2_u0_n93 ) );
  NAND2_X1 u1_u2_u0_U46 (.ZN( u1_u2_u0_n112 ) , .A2( u1_u2_u0_n92 ) , .A1( u1_u2_u0_n93 ) );
  OR3_X1 u1_u2_u0_U47 (.A3( u1_u2_u0_n152 ) , .A2( u1_u2_u0_n153 ) , .A1( u1_u2_u0_n154 ) , .ZN( u1_u2_u0_n155 ) );
  AOI21_X1 u1_u2_u0_U48 (.B2( u1_u2_u0_n150 ) , .B1( u1_u2_u0_n151 ) , .ZN( u1_u2_u0_n152 ) , .A( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U49 (.A( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n145 ) , .B1( u1_u2_u0_n146 ) , .ZN( u1_u2_u0_n154 ) );
  AOI21_X1 u1_u2_u0_U5 (.B2( u1_u2_u0_n131 ) , .ZN( u1_u2_u0_n134 ) , .B1( u1_u2_u0_n151 ) , .A( u1_u2_u0_n158 ) );
  AOI21_X1 u1_u2_u0_U50 (.A( u1_u2_u0_n147 ) , .B2( u1_u2_u0_n148 ) , .B1( u1_u2_u0_n149 ) , .ZN( u1_u2_u0_n153 ) );
  INV_X1 u1_u2_u0_U51 (.ZN( u1_u2_u0_n171 ) , .A( u1_u2_u0_n99 ) );
  OAI211_X1 u1_u2_u0_U52 (.C2( u1_u2_u0_n140 ) , .C1( u1_u2_u0_n161 ) , .A( u1_u2_u0_n169 ) , .B( u1_u2_u0_n98 ) , .ZN( u1_u2_u0_n99 ) );
  AOI211_X1 u1_u2_u0_U53 (.C1( u1_u2_u0_n118 ) , .A( u1_u2_u0_n123 ) , .B( u1_u2_u0_n96 ) , .C2( u1_u2_u0_n97 ) , .ZN( u1_u2_u0_n98 ) );
  INV_X1 u1_u2_u0_U54 (.ZN( u1_u2_u0_n169 ) , .A( u1_u2_u0_n91 ) );
  NOR2_X1 u1_u2_u0_U55 (.A2( u1_u2_X_6 ) , .ZN( u1_u2_u0_n100 ) , .A1( u1_u2_u0_n162 ) );
  NOR2_X1 u1_u2_u0_U56 (.A2( u1_u2_X_4 ) , .A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n118 ) );
  NOR2_X1 u1_u2_u0_U57 (.A2( u1_u2_X_2 ) , .ZN( u1_u2_u0_n103 ) , .A1( u1_u2_u0_n164 ) );
  NOR2_X1 u1_u2_u0_U58 (.A2( u1_u2_X_1 ) , .A1( u1_u2_X_2 ) , .ZN( u1_u2_u0_n92 ) );
  NOR2_X1 u1_u2_u0_U59 (.A2( u1_u2_X_1 ) , .ZN( u1_u2_u0_n101 ) , .A1( u1_u2_u0_n163 ) );
  NOR2_X1 u1_u2_u0_U6 (.A1( u1_u2_u0_n108 ) , .ZN( u1_u2_u0_n123 ) , .A2( u1_u2_u0_n158 ) );
  NAND2_X1 u1_u2_u0_U60 (.A2( u1_u2_X_4 ) , .A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n144 ) );
  NOR2_X1 u1_u2_u0_U61 (.A2( u1_u2_X_5 ) , .ZN( u1_u2_u0_n136 ) , .A1( u1_u2_u0_n159 ) );
  NAND2_X1 u1_u2_u0_U62 (.A1( u1_u2_X_5 ) , .ZN( u1_u2_u0_n138 ) , .A2( u1_u2_u0_n159 ) );
  AND2_X1 u1_u2_u0_U63 (.A2( u1_u2_X_3 ) , .A1( u1_u2_X_6 ) , .ZN( u1_u2_u0_n102 ) );
  AND2_X1 u1_u2_u0_U64 (.A1( u1_u2_X_6 ) , .A2( u1_u2_u0_n162 ) , .ZN( u1_u2_u0_n93 ) );
  INV_X1 u1_u2_u0_U65 (.A( u1_u2_X_4 ) , .ZN( u1_u2_u0_n159 ) );
  INV_X1 u1_u2_u0_U66 (.A( u1_u2_X_1 ) , .ZN( u1_u2_u0_n164 ) );
  INV_X1 u1_u2_u0_U67 (.A( u1_u2_X_2 ) , .ZN( u1_u2_u0_n163 ) );
  INV_X1 u1_u2_u0_U68 (.ZN( u1_u2_u0_n174 ) , .A( u1_u2_u0_n89 ) );
  AOI211_X1 u1_u2_u0_U69 (.B( u1_u2_u0_n104 ) , .A( u1_u2_u0_n105 ) , .ZN( u1_u2_u0_n106 ) , .C2( u1_u2_u0_n113 ) , .C1( u1_u2_u0_n160 ) );
  OAI21_X1 u1_u2_u0_U7 (.B1( u1_u2_u0_n150 ) , .B2( u1_u2_u0_n158 ) , .A( u1_u2_u0_n172 ) , .ZN( u1_u2_u0_n89 ) );
  OR4_X1 u1_u2_u0_U70 (.ZN( u1_out2_17 ) , .A4( u1_u2_u0_n122 ) , .A2( u1_u2_u0_n123 ) , .A1( u1_u2_u0_n124 ) , .A3( u1_u2_u0_n170 ) );
  AOI21_X1 u1_u2_u0_U71 (.B2( u1_u2_u0_n107 ) , .ZN( u1_u2_u0_n124 ) , .B1( u1_u2_u0_n128 ) , .A( u1_u2_u0_n161 ) );
  INV_X1 u1_u2_u0_U72 (.A( u1_u2_u0_n111 ) , .ZN( u1_u2_u0_n170 ) );
  OR4_X1 u1_u2_u0_U73 (.ZN( u1_out2_31 ) , .A4( u1_u2_u0_n155 ) , .A2( u1_u2_u0_n156 ) , .A1( u1_u2_u0_n157 ) , .A3( u1_u2_u0_n173 ) );
  AOI21_X1 u1_u2_u0_U74 (.A( u1_u2_u0_n138 ) , .B2( u1_u2_u0_n139 ) , .B1( u1_u2_u0_n140 ) , .ZN( u1_u2_u0_n157 ) );
  AOI21_X1 u1_u2_u0_U75 (.B2( u1_u2_u0_n141 ) , .B1( u1_u2_u0_n142 ) , .ZN( u1_u2_u0_n156 ) , .A( u1_u2_u0_n161 ) );
  INV_X1 u1_u2_u0_U76 (.A( u1_u2_u0_n126 ) , .ZN( u1_u2_u0_n168 ) );
  AOI211_X1 u1_u2_u0_U77 (.B( u1_u2_u0_n133 ) , .A( u1_u2_u0_n134 ) , .C2( u1_u2_u0_n135 ) , .C1( u1_u2_u0_n136 ) , .ZN( u1_u2_u0_n137 ) );
  AOI21_X1 u1_u2_u0_U78 (.B1( u1_u2_u0_n132 ) , .ZN( u1_u2_u0_n133 ) , .A( u1_u2_u0_n144 ) , .B2( u1_u2_u0_n166 ) );
  OAI22_X1 u1_u2_u0_U79 (.ZN( u1_u2_u0_n105 ) , .A2( u1_u2_u0_n132 ) , .B1( u1_u2_u0_n146 ) , .A1( u1_u2_u0_n147 ) , .B2( u1_u2_u0_n161 ) );
  AND2_X1 u1_u2_u0_U8 (.A1( u1_u2_u0_n114 ) , .A2( u1_u2_u0_n121 ) , .ZN( u1_u2_u0_n146 ) );
  NAND2_X1 u1_u2_u0_U80 (.ZN( u1_u2_u0_n110 ) , .A2( u1_u2_u0_n132 ) , .A1( u1_u2_u0_n145 ) );
  INV_X1 u1_u2_u0_U81 (.A( u1_u2_u0_n119 ) , .ZN( u1_u2_u0_n167 ) );
  NAND2_X1 u1_u2_u0_U82 (.A2( u1_u2_u0_n103 ) , .ZN( u1_u2_u0_n140 ) , .A1( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U83 (.A1( u1_u2_u0_n101 ) , .ZN( u1_u2_u0_n130 ) , .A2( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U84 (.ZN( u1_u2_u0_n108 ) , .A1( u1_u2_u0_n92 ) , .A2( u1_u2_u0_n94 ) );
  NAND2_X1 u1_u2_u0_U85 (.ZN( u1_u2_u0_n142 ) , .A1( u1_u2_u0_n94 ) , .A2( u1_u2_u0_n95 ) );
  INV_X1 u1_u2_u0_U86 (.A( u1_u2_X_3 ) , .ZN( u1_u2_u0_n162 ) );
  NOR2_X1 u1_u2_u0_U87 (.A2( u1_u2_X_3 ) , .A1( u1_u2_X_6 ) , .ZN( u1_u2_u0_n94 ) );
  NAND3_X1 u1_u2_u0_U88 (.ZN( u1_out2_23 ) , .A3( u1_u2_u0_n137 ) , .A1( u1_u2_u0_n168 ) , .A2( u1_u2_u0_n171 ) );
  NAND3_X1 u1_u2_u0_U89 (.A3( u1_u2_u0_n127 ) , .A2( u1_u2_u0_n128 ) , .ZN( u1_u2_u0_n135 ) , .A1( u1_u2_u0_n150 ) );
  AND2_X1 u1_u2_u0_U9 (.A1( u1_u2_u0_n131 ) , .ZN( u1_u2_u0_n141 ) , .A2( u1_u2_u0_n150 ) );
  NAND3_X1 u1_u2_u0_U90 (.ZN( u1_u2_u0_n117 ) , .A3( u1_u2_u0_n132 ) , .A2( u1_u2_u0_n139 ) , .A1( u1_u2_u0_n148 ) );
  NAND3_X1 u1_u2_u0_U91 (.ZN( u1_u2_u0_n109 ) , .A2( u1_u2_u0_n114 ) , .A3( u1_u2_u0_n140 ) , .A1( u1_u2_u0_n149 ) );
  NAND3_X1 u1_u2_u0_U92 (.ZN( u1_out2_9 ) , .A3( u1_u2_u0_n106 ) , .A2( u1_u2_u0_n171 ) , .A1( u1_u2_u0_n174 ) );
  NAND3_X1 u1_u2_u0_U93 (.A2( u1_u2_u0_n128 ) , .A1( u1_u2_u0_n132 ) , .A3( u1_u2_u0_n146 ) , .ZN( u1_u2_u0_n97 ) );
  NOR2_X1 u1_u2_u1_U10 (.A1( u1_u2_u1_n112 ) , .A2( u1_u2_u1_n116 ) , .ZN( u1_u2_u1_n118 ) );
  NAND3_X1 u1_u2_u1_U100 (.ZN( u1_u2_u1_n113 ) , .A1( u1_u2_u1_n120 ) , .A3( u1_u2_u1_n133 ) , .A2( u1_u2_u1_n155 ) );
  OAI21_X1 u1_u2_u1_U11 (.ZN( u1_u2_u1_n101 ) , .B1( u1_u2_u1_n141 ) , .A( u1_u2_u1_n146 ) , .B2( u1_u2_u1_n183 ) );
  AOI21_X1 u1_u2_u1_U12 (.B2( u1_u2_u1_n155 ) , .B1( u1_u2_u1_n156 ) , .ZN( u1_u2_u1_n157 ) , .A( u1_u2_u1_n174 ) );
  OR4_X1 u1_u2_u1_U13 (.A4( u1_u2_u1_n106 ) , .A3( u1_u2_u1_n107 ) , .ZN( u1_u2_u1_n108 ) , .A1( u1_u2_u1_n117 ) , .A2( u1_u2_u1_n184 ) );
  AOI21_X1 u1_u2_u1_U14 (.ZN( u1_u2_u1_n106 ) , .A( u1_u2_u1_n112 ) , .B1( u1_u2_u1_n154 ) , .B2( u1_u2_u1_n156 ) );
  INV_X1 u1_u2_u1_U15 (.A( u1_u2_u1_n101 ) , .ZN( u1_u2_u1_n184 ) );
  AOI21_X1 u1_u2_u1_U16 (.ZN( u1_u2_u1_n107 ) , .B1( u1_u2_u1_n134 ) , .B2( u1_u2_u1_n149 ) , .A( u1_u2_u1_n174 ) );
  NAND2_X1 u1_u2_u1_U17 (.ZN( u1_u2_u1_n140 ) , .A2( u1_u2_u1_n150 ) , .A1( u1_u2_u1_n155 ) );
  NAND2_X1 u1_u2_u1_U18 (.A1( u1_u2_u1_n131 ) , .ZN( u1_u2_u1_n147 ) , .A2( u1_u2_u1_n153 ) );
  INV_X1 u1_u2_u1_U19 (.A( u1_u2_u1_n139 ) , .ZN( u1_u2_u1_n174 ) );
  INV_X1 u1_u2_u1_U20 (.A( u1_u2_u1_n112 ) , .ZN( u1_u2_u1_n171 ) );
  NAND2_X1 u1_u2_u1_U21 (.ZN( u1_u2_u1_n141 ) , .A1( u1_u2_u1_n153 ) , .A2( u1_u2_u1_n156 ) );
  AND2_X1 u1_u2_u1_U22 (.A1( u1_u2_u1_n123 ) , .ZN( u1_u2_u1_n134 ) , .A2( u1_u2_u1_n161 ) );
  NAND2_X1 u1_u2_u1_U23 (.A2( u1_u2_u1_n115 ) , .A1( u1_u2_u1_n116 ) , .ZN( u1_u2_u1_n148 ) );
  NAND2_X1 u1_u2_u1_U24 (.A2( u1_u2_u1_n133 ) , .A1( u1_u2_u1_n135 ) , .ZN( u1_u2_u1_n159 ) );
  NAND2_X1 u1_u2_u1_U25 (.A2( u1_u2_u1_n115 ) , .A1( u1_u2_u1_n120 ) , .ZN( u1_u2_u1_n132 ) );
  INV_X1 u1_u2_u1_U26 (.A( u1_u2_u1_n154 ) , .ZN( u1_u2_u1_n178 ) );
  INV_X1 u1_u2_u1_U27 (.A( u1_u2_u1_n151 ) , .ZN( u1_u2_u1_n183 ) );
  AND2_X1 u1_u2_u1_U28 (.A1( u1_u2_u1_n129 ) , .A2( u1_u2_u1_n133 ) , .ZN( u1_u2_u1_n149 ) );
  INV_X1 u1_u2_u1_U29 (.A( u1_u2_u1_n131 ) , .ZN( u1_u2_u1_n180 ) );
  INV_X1 u1_u2_u1_U3 (.A( u1_u2_u1_n159 ) , .ZN( u1_u2_u1_n182 ) );
  OAI221_X1 u1_u2_u1_U30 (.A( u1_u2_u1_n119 ) , .C2( u1_u2_u1_n129 ) , .ZN( u1_u2_u1_n138 ) , .B2( u1_u2_u1_n152 ) , .C1( u1_u2_u1_n174 ) , .B1( u1_u2_u1_n187 ) );
  INV_X1 u1_u2_u1_U31 (.A( u1_u2_u1_n148 ) , .ZN( u1_u2_u1_n187 ) );
  AOI211_X1 u1_u2_u1_U32 (.B( u1_u2_u1_n117 ) , .A( u1_u2_u1_n118 ) , .ZN( u1_u2_u1_n119 ) , .C2( u1_u2_u1_n146 ) , .C1( u1_u2_u1_n159 ) );
  NOR2_X1 u1_u2_u1_U33 (.A1( u1_u2_u1_n168 ) , .A2( u1_u2_u1_n176 ) , .ZN( u1_u2_u1_n98 ) );
  AOI211_X1 u1_u2_u1_U34 (.B( u1_u2_u1_n162 ) , .A( u1_u2_u1_n163 ) , .C2( u1_u2_u1_n164 ) , .ZN( u1_u2_u1_n165 ) , .C1( u1_u2_u1_n171 ) );
  AOI21_X1 u1_u2_u1_U35 (.A( u1_u2_u1_n160 ) , .B2( u1_u2_u1_n161 ) , .ZN( u1_u2_u1_n162 ) , .B1( u1_u2_u1_n182 ) );
  OR2_X1 u1_u2_u1_U36 (.A2( u1_u2_u1_n157 ) , .A1( u1_u2_u1_n158 ) , .ZN( u1_u2_u1_n163 ) );
  OAI21_X1 u1_u2_u1_U37 (.B2( u1_u2_u1_n123 ) , .ZN( u1_u2_u1_n145 ) , .B1( u1_u2_u1_n160 ) , .A( u1_u2_u1_n185 ) );
  INV_X1 u1_u2_u1_U38 (.A( u1_u2_u1_n122 ) , .ZN( u1_u2_u1_n185 ) );
  AOI21_X1 u1_u2_u1_U39 (.B2( u1_u2_u1_n120 ) , .B1( u1_u2_u1_n121 ) , .ZN( u1_u2_u1_n122 ) , .A( u1_u2_u1_n128 ) );
  AOI221_X1 u1_u2_u1_U4 (.A( u1_u2_u1_n138 ) , .C2( u1_u2_u1_n139 ) , .C1( u1_u2_u1_n140 ) , .B2( u1_u2_u1_n141 ) , .ZN( u1_u2_u1_n142 ) , .B1( u1_u2_u1_n175 ) );
  NAND2_X1 u1_u2_u1_U40 (.A1( u1_u2_u1_n128 ) , .ZN( u1_u2_u1_n146 ) , .A2( u1_u2_u1_n160 ) );
  NAND2_X1 u1_u2_u1_U41 (.A2( u1_u2_u1_n112 ) , .ZN( u1_u2_u1_n139 ) , .A1( u1_u2_u1_n152 ) );
  NAND2_X1 u1_u2_u1_U42 (.A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n156 ) , .A2( u1_u2_u1_n99 ) );
  AOI221_X1 u1_u2_u1_U43 (.B1( u1_u2_u1_n140 ) , .ZN( u1_u2_u1_n167 ) , .B2( u1_u2_u1_n172 ) , .C2( u1_u2_u1_n175 ) , .C1( u1_u2_u1_n178 ) , .A( u1_u2_u1_n188 ) );
  INV_X1 u1_u2_u1_U44 (.ZN( u1_u2_u1_n188 ) , .A( u1_u2_u1_n97 ) );
  AOI211_X1 u1_u2_u1_U45 (.A( u1_u2_u1_n118 ) , .C1( u1_u2_u1_n132 ) , .C2( u1_u2_u1_n139 ) , .B( u1_u2_u1_n96 ) , .ZN( u1_u2_u1_n97 ) );
  AOI21_X1 u1_u2_u1_U46 (.B2( u1_u2_u1_n121 ) , .B1( u1_u2_u1_n135 ) , .A( u1_u2_u1_n152 ) , .ZN( u1_u2_u1_n96 ) );
  NOR2_X1 u1_u2_u1_U47 (.ZN( u1_u2_u1_n117 ) , .A1( u1_u2_u1_n121 ) , .A2( u1_u2_u1_n160 ) );
  AOI21_X1 u1_u2_u1_U48 (.A( u1_u2_u1_n128 ) , .B2( u1_u2_u1_n129 ) , .ZN( u1_u2_u1_n130 ) , .B1( u1_u2_u1_n150 ) );
  NAND2_X1 u1_u2_u1_U49 (.ZN( u1_u2_u1_n112 ) , .A1( u1_u2_u1_n169 ) , .A2( u1_u2_u1_n170 ) );
  AOI211_X1 u1_u2_u1_U5 (.ZN( u1_u2_u1_n124 ) , .A( u1_u2_u1_n138 ) , .C2( u1_u2_u1_n139 ) , .B( u1_u2_u1_n145 ) , .C1( u1_u2_u1_n147 ) );
  NAND2_X1 u1_u2_u1_U50 (.ZN( u1_u2_u1_n129 ) , .A2( u1_u2_u1_n95 ) , .A1( u1_u2_u1_n98 ) );
  NAND2_X1 u1_u2_u1_U51 (.A1( u1_u2_u1_n102 ) , .ZN( u1_u2_u1_n154 ) , .A2( u1_u2_u1_n99 ) );
  NAND2_X1 u1_u2_u1_U52 (.A2( u1_u2_u1_n100 ) , .ZN( u1_u2_u1_n135 ) , .A1( u1_u2_u1_n99 ) );
  AOI21_X1 u1_u2_u1_U53 (.A( u1_u2_u1_n152 ) , .B2( u1_u2_u1_n153 ) , .B1( u1_u2_u1_n154 ) , .ZN( u1_u2_u1_n158 ) );
  INV_X1 u1_u2_u1_U54 (.A( u1_u2_u1_n160 ) , .ZN( u1_u2_u1_n175 ) );
  NAND2_X1 u1_u2_u1_U55 (.A1( u1_u2_u1_n100 ) , .ZN( u1_u2_u1_n116 ) , .A2( u1_u2_u1_n95 ) );
  NAND2_X1 u1_u2_u1_U56 (.A1( u1_u2_u1_n102 ) , .ZN( u1_u2_u1_n131 ) , .A2( u1_u2_u1_n95 ) );
  NAND2_X1 u1_u2_u1_U57 (.A2( u1_u2_u1_n104 ) , .ZN( u1_u2_u1_n121 ) , .A1( u1_u2_u1_n98 ) );
  NAND2_X1 u1_u2_u1_U58 (.A1( u1_u2_u1_n103 ) , .ZN( u1_u2_u1_n153 ) , .A2( u1_u2_u1_n98 ) );
  NAND2_X1 u1_u2_u1_U59 (.A2( u1_u2_u1_n104 ) , .A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n133 ) );
  AOI22_X1 u1_u2_u1_U6 (.B2( u1_u2_u1_n113 ) , .A2( u1_u2_u1_n114 ) , .ZN( u1_u2_u1_n125 ) , .A1( u1_u2_u1_n171 ) , .B1( u1_u2_u1_n173 ) );
  NAND2_X1 u1_u2_u1_U60 (.ZN( u1_u2_u1_n150 ) , .A2( u1_u2_u1_n98 ) , .A1( u1_u2_u1_n99 ) );
  NAND2_X1 u1_u2_u1_U61 (.A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n155 ) , .A2( u1_u2_u1_n95 ) );
  OAI21_X1 u1_u2_u1_U62 (.ZN( u1_u2_u1_n109 ) , .B1( u1_u2_u1_n129 ) , .B2( u1_u2_u1_n160 ) , .A( u1_u2_u1_n167 ) );
  NAND2_X1 u1_u2_u1_U63 (.A2( u1_u2_u1_n100 ) , .A1( u1_u2_u1_n103 ) , .ZN( u1_u2_u1_n120 ) );
  NAND2_X1 u1_u2_u1_U64 (.A1( u1_u2_u1_n102 ) , .A2( u1_u2_u1_n104 ) , .ZN( u1_u2_u1_n115 ) );
  NAND2_X1 u1_u2_u1_U65 (.A2( u1_u2_u1_n100 ) , .A1( u1_u2_u1_n104 ) , .ZN( u1_u2_u1_n151 ) );
  NAND2_X1 u1_u2_u1_U66 (.A2( u1_u2_u1_n103 ) , .A1( u1_u2_u1_n105 ) , .ZN( u1_u2_u1_n161 ) );
  INV_X1 u1_u2_u1_U67 (.A( u1_u2_u1_n152 ) , .ZN( u1_u2_u1_n173 ) );
  INV_X1 u1_u2_u1_U68 (.A( u1_u2_u1_n128 ) , .ZN( u1_u2_u1_n172 ) );
  NAND2_X1 u1_u2_u1_U69 (.A2( u1_u2_u1_n102 ) , .A1( u1_u2_u1_n103 ) , .ZN( u1_u2_u1_n123 ) );
  NAND2_X1 u1_u2_u1_U7 (.ZN( u1_u2_u1_n114 ) , .A1( u1_u2_u1_n134 ) , .A2( u1_u2_u1_n156 ) );
  NOR2_X1 u1_u2_u1_U70 (.A2( u1_u2_X_7 ) , .A1( u1_u2_X_8 ) , .ZN( u1_u2_u1_n95 ) );
  NOR2_X1 u1_u2_u1_U71 (.A1( u1_u2_X_12 ) , .A2( u1_u2_X_9 ) , .ZN( u1_u2_u1_n100 ) );
  NOR2_X1 u1_u2_u1_U72 (.A2( u1_u2_X_8 ) , .A1( u1_u2_u1_n177 ) , .ZN( u1_u2_u1_n99 ) );
  NOR2_X1 u1_u2_u1_U73 (.A2( u1_u2_X_12 ) , .ZN( u1_u2_u1_n102 ) , .A1( u1_u2_u1_n176 ) );
  NOR2_X1 u1_u2_u1_U74 (.A2( u1_u2_X_9 ) , .ZN( u1_u2_u1_n105 ) , .A1( u1_u2_u1_n168 ) );
  NAND2_X1 u1_u2_u1_U75 (.A1( u1_u2_X_10 ) , .ZN( u1_u2_u1_n160 ) , .A2( u1_u2_u1_n169 ) );
  NAND2_X1 u1_u2_u1_U76 (.A2( u1_u2_X_10 ) , .A1( u1_u2_X_11 ) , .ZN( u1_u2_u1_n152 ) );
  NAND2_X1 u1_u2_u1_U77 (.A1( u1_u2_X_11 ) , .ZN( u1_u2_u1_n128 ) , .A2( u1_u2_u1_n170 ) );
  AND2_X1 u1_u2_u1_U78 (.A2( u1_u2_X_7 ) , .A1( u1_u2_X_8 ) , .ZN( u1_u2_u1_n104 ) );
  AND2_X1 u1_u2_u1_U79 (.A1( u1_u2_X_8 ) , .ZN( u1_u2_u1_n103 ) , .A2( u1_u2_u1_n177 ) );
  AOI22_X1 u1_u2_u1_U8 (.B2( u1_u2_u1_n136 ) , .A2( u1_u2_u1_n137 ) , .ZN( u1_u2_u1_n143 ) , .A1( u1_u2_u1_n171 ) , .B1( u1_u2_u1_n173 ) );
  INV_X1 u1_u2_u1_U80 (.A( u1_u2_X_10 ) , .ZN( u1_u2_u1_n170 ) );
  INV_X1 u1_u2_u1_U81 (.A( u1_u2_X_9 ) , .ZN( u1_u2_u1_n176 ) );
  INV_X1 u1_u2_u1_U82 (.A( u1_u2_X_11 ) , .ZN( u1_u2_u1_n169 ) );
  INV_X1 u1_u2_u1_U83 (.A( u1_u2_X_12 ) , .ZN( u1_u2_u1_n168 ) );
  INV_X1 u1_u2_u1_U84 (.A( u1_u2_X_7 ) , .ZN( u1_u2_u1_n177 ) );
  NAND4_X1 u1_u2_u1_U85 (.ZN( u1_out2_18 ) , .A4( u1_u2_u1_n165 ) , .A3( u1_u2_u1_n166 ) , .A1( u1_u2_u1_n167 ) , .A2( u1_u2_u1_n186 ) );
  AOI22_X1 u1_u2_u1_U86 (.B2( u1_u2_u1_n146 ) , .B1( u1_u2_u1_n147 ) , .A2( u1_u2_u1_n148 ) , .ZN( u1_u2_u1_n166 ) , .A1( u1_u2_u1_n172 ) );
  INV_X1 u1_u2_u1_U87 (.A( u1_u2_u1_n145 ) , .ZN( u1_u2_u1_n186 ) );
  NAND4_X1 u1_u2_u1_U88 (.ZN( u1_out2_2 ) , .A4( u1_u2_u1_n142 ) , .A3( u1_u2_u1_n143 ) , .A2( u1_u2_u1_n144 ) , .A1( u1_u2_u1_n179 ) );
  OAI21_X1 u1_u2_u1_U89 (.B2( u1_u2_u1_n132 ) , .ZN( u1_u2_u1_n144 ) , .A( u1_u2_u1_n146 ) , .B1( u1_u2_u1_n180 ) );
  INV_X1 u1_u2_u1_U9 (.A( u1_u2_u1_n147 ) , .ZN( u1_u2_u1_n181 ) );
  INV_X1 u1_u2_u1_U90 (.A( u1_u2_u1_n130 ) , .ZN( u1_u2_u1_n179 ) );
  NAND4_X1 u1_u2_u1_U91 (.ZN( u1_out2_28 ) , .A4( u1_u2_u1_n124 ) , .A3( u1_u2_u1_n125 ) , .A2( u1_u2_u1_n126 ) , .A1( u1_u2_u1_n127 ) );
  OAI21_X1 u1_u2_u1_U92 (.ZN( u1_u2_u1_n127 ) , .B2( u1_u2_u1_n139 ) , .B1( u1_u2_u1_n175 ) , .A( u1_u2_u1_n183 ) );
  OAI21_X1 u1_u2_u1_U93 (.ZN( u1_u2_u1_n126 ) , .B2( u1_u2_u1_n140 ) , .A( u1_u2_u1_n146 ) , .B1( u1_u2_u1_n178 ) );
  OR4_X1 u1_u2_u1_U94 (.ZN( u1_out2_13 ) , .A4( u1_u2_u1_n108 ) , .A3( u1_u2_u1_n109 ) , .A2( u1_u2_u1_n110 ) , .A1( u1_u2_u1_n111 ) );
  AOI21_X1 u1_u2_u1_U95 (.ZN( u1_u2_u1_n111 ) , .A( u1_u2_u1_n128 ) , .B2( u1_u2_u1_n131 ) , .B1( u1_u2_u1_n135 ) );
  AOI21_X1 u1_u2_u1_U96 (.ZN( u1_u2_u1_n110 ) , .A( u1_u2_u1_n116 ) , .B1( u1_u2_u1_n152 ) , .B2( u1_u2_u1_n160 ) );
  NAND3_X1 u1_u2_u1_U97 (.A3( u1_u2_u1_n149 ) , .A2( u1_u2_u1_n150 ) , .A1( u1_u2_u1_n151 ) , .ZN( u1_u2_u1_n164 ) );
  NAND3_X1 u1_u2_u1_U98 (.A3( u1_u2_u1_n134 ) , .A2( u1_u2_u1_n135 ) , .ZN( u1_u2_u1_n136 ) , .A1( u1_u2_u1_n151 ) );
  NAND3_X1 u1_u2_u1_U99 (.A1( u1_u2_u1_n133 ) , .ZN( u1_u2_u1_n137 ) , .A2( u1_u2_u1_n154 ) , .A3( u1_u2_u1_n181 ) );
  OAI22_X1 u1_u2_u2_U10 (.B1( u1_u2_u2_n151 ) , .A2( u1_u2_u2_n152 ) , .A1( u1_u2_u2_n153 ) , .ZN( u1_u2_u2_n160 ) , .B2( u1_u2_u2_n168 ) );
  NAND3_X1 u1_u2_u2_U100 (.A2( u1_u2_u2_n100 ) , .A1( u1_u2_u2_n104 ) , .A3( u1_u2_u2_n138 ) , .ZN( u1_u2_u2_n98 ) );
  NOR3_X1 u1_u2_u2_U11 (.A1( u1_u2_u2_n150 ) , .ZN( u1_u2_u2_n151 ) , .A3( u1_u2_u2_n175 ) , .A2( u1_u2_u2_n188 ) );
  AOI21_X1 u1_u2_u2_U12 (.B2( u1_u2_u2_n123 ) , .ZN( u1_u2_u2_n125 ) , .A( u1_u2_u2_n171 ) , .B1( u1_u2_u2_n184 ) );
  INV_X1 u1_u2_u2_U13 (.A( u1_u2_u2_n150 ) , .ZN( u1_u2_u2_n184 ) );
  AOI21_X1 u1_u2_u2_U14 (.ZN( u1_u2_u2_n144 ) , .B2( u1_u2_u2_n155 ) , .A( u1_u2_u2_n172 ) , .B1( u1_u2_u2_n185 ) );
  AOI21_X1 u1_u2_u2_U15 (.B2( u1_u2_u2_n143 ) , .ZN( u1_u2_u2_n145 ) , .B1( u1_u2_u2_n152 ) , .A( u1_u2_u2_n171 ) );
  INV_X1 u1_u2_u2_U16 (.A( u1_u2_u2_n156 ) , .ZN( u1_u2_u2_n171 ) );
  INV_X1 u1_u2_u2_U17 (.A( u1_u2_u2_n120 ) , .ZN( u1_u2_u2_n188 ) );
  NAND2_X1 u1_u2_u2_U18 (.A2( u1_u2_u2_n122 ) , .ZN( u1_u2_u2_n150 ) , .A1( u1_u2_u2_n152 ) );
  INV_X1 u1_u2_u2_U19 (.A( u1_u2_u2_n153 ) , .ZN( u1_u2_u2_n170 ) );
  INV_X1 u1_u2_u2_U20 (.A( u1_u2_u2_n137 ) , .ZN( u1_u2_u2_n173 ) );
  NAND2_X1 u1_u2_u2_U21 (.A1( u1_u2_u2_n132 ) , .A2( u1_u2_u2_n139 ) , .ZN( u1_u2_u2_n157 ) );
  INV_X1 u1_u2_u2_U22 (.A( u1_u2_u2_n113 ) , .ZN( u1_u2_u2_n178 ) );
  INV_X1 u1_u2_u2_U23 (.A( u1_u2_u2_n139 ) , .ZN( u1_u2_u2_n175 ) );
  INV_X1 u1_u2_u2_U24 (.A( u1_u2_u2_n155 ) , .ZN( u1_u2_u2_n181 ) );
  INV_X1 u1_u2_u2_U25 (.A( u1_u2_u2_n119 ) , .ZN( u1_u2_u2_n177 ) );
  INV_X1 u1_u2_u2_U26 (.A( u1_u2_u2_n116 ) , .ZN( u1_u2_u2_n180 ) );
  INV_X1 u1_u2_u2_U27 (.A( u1_u2_u2_n131 ) , .ZN( u1_u2_u2_n179 ) );
  INV_X1 u1_u2_u2_U28 (.A( u1_u2_u2_n154 ) , .ZN( u1_u2_u2_n176 ) );
  NAND2_X1 u1_u2_u2_U29 (.A2( u1_u2_u2_n116 ) , .A1( u1_u2_u2_n117 ) , .ZN( u1_u2_u2_n118 ) );
  NOR2_X1 u1_u2_u2_U3 (.ZN( u1_u2_u2_n121 ) , .A2( u1_u2_u2_n177 ) , .A1( u1_u2_u2_n180 ) );
  INV_X1 u1_u2_u2_U30 (.A( u1_u2_u2_n132 ) , .ZN( u1_u2_u2_n182 ) );
  INV_X1 u1_u2_u2_U31 (.A( u1_u2_u2_n158 ) , .ZN( u1_u2_u2_n183 ) );
  OAI21_X1 u1_u2_u2_U32 (.A( u1_u2_u2_n156 ) , .B1( u1_u2_u2_n157 ) , .ZN( u1_u2_u2_n158 ) , .B2( u1_u2_u2_n179 ) );
  NOR2_X1 u1_u2_u2_U33 (.ZN( u1_u2_u2_n156 ) , .A1( u1_u2_u2_n166 ) , .A2( u1_u2_u2_n169 ) );
  NOR2_X1 u1_u2_u2_U34 (.A2( u1_u2_u2_n114 ) , .ZN( u1_u2_u2_n137 ) , .A1( u1_u2_u2_n140 ) );
  NOR2_X1 u1_u2_u2_U35 (.A2( u1_u2_u2_n138 ) , .ZN( u1_u2_u2_n153 ) , .A1( u1_u2_u2_n156 ) );
  AOI211_X1 u1_u2_u2_U36 (.ZN( u1_u2_u2_n130 ) , .C1( u1_u2_u2_n138 ) , .C2( u1_u2_u2_n179 ) , .B( u1_u2_u2_n96 ) , .A( u1_u2_u2_n97 ) );
  OAI22_X1 u1_u2_u2_U37 (.B1( u1_u2_u2_n133 ) , .A2( u1_u2_u2_n137 ) , .A1( u1_u2_u2_n152 ) , .B2( u1_u2_u2_n168 ) , .ZN( u1_u2_u2_n97 ) );
  OAI221_X1 u1_u2_u2_U38 (.B1( u1_u2_u2_n113 ) , .C1( u1_u2_u2_n132 ) , .A( u1_u2_u2_n149 ) , .B2( u1_u2_u2_n171 ) , .C2( u1_u2_u2_n172 ) , .ZN( u1_u2_u2_n96 ) );
  OAI221_X1 u1_u2_u2_U39 (.A( u1_u2_u2_n115 ) , .C2( u1_u2_u2_n123 ) , .B2( u1_u2_u2_n143 ) , .B1( u1_u2_u2_n153 ) , .ZN( u1_u2_u2_n163 ) , .C1( u1_u2_u2_n168 ) );
  INV_X1 u1_u2_u2_U4 (.A( u1_u2_u2_n134 ) , .ZN( u1_u2_u2_n185 ) );
  OAI21_X1 u1_u2_u2_U40 (.A( u1_u2_u2_n114 ) , .ZN( u1_u2_u2_n115 ) , .B1( u1_u2_u2_n176 ) , .B2( u1_u2_u2_n178 ) );
  OAI221_X1 u1_u2_u2_U41 (.A( u1_u2_u2_n135 ) , .B2( u1_u2_u2_n136 ) , .B1( u1_u2_u2_n137 ) , .ZN( u1_u2_u2_n162 ) , .C2( u1_u2_u2_n167 ) , .C1( u1_u2_u2_n185 ) );
  AND3_X1 u1_u2_u2_U42 (.A3( u1_u2_u2_n131 ) , .A2( u1_u2_u2_n132 ) , .A1( u1_u2_u2_n133 ) , .ZN( u1_u2_u2_n136 ) );
  AOI22_X1 u1_u2_u2_U43 (.ZN( u1_u2_u2_n135 ) , .B1( u1_u2_u2_n140 ) , .A1( u1_u2_u2_n156 ) , .B2( u1_u2_u2_n180 ) , .A2( u1_u2_u2_n188 ) );
  AOI21_X1 u1_u2_u2_U44 (.ZN( u1_u2_u2_n149 ) , .B1( u1_u2_u2_n173 ) , .B2( u1_u2_u2_n188 ) , .A( u1_u2_u2_n95 ) );
  AND3_X1 u1_u2_u2_U45 (.A2( u1_u2_u2_n100 ) , .A1( u1_u2_u2_n104 ) , .A3( u1_u2_u2_n156 ) , .ZN( u1_u2_u2_n95 ) );
  OAI21_X1 u1_u2_u2_U46 (.A( u1_u2_u2_n101 ) , .B2( u1_u2_u2_n121 ) , .B1( u1_u2_u2_n153 ) , .ZN( u1_u2_u2_n164 ) );
  NAND2_X1 u1_u2_u2_U47 (.A2( u1_u2_u2_n100 ) , .A1( u1_u2_u2_n107 ) , .ZN( u1_u2_u2_n155 ) );
  NAND2_X1 u1_u2_u2_U48 (.A2( u1_u2_u2_n105 ) , .A1( u1_u2_u2_n108 ) , .ZN( u1_u2_u2_n143 ) );
  NAND2_X1 u1_u2_u2_U49 (.A1( u1_u2_u2_n104 ) , .A2( u1_u2_u2_n106 ) , .ZN( u1_u2_u2_n152 ) );
  NOR4_X1 u1_u2_u2_U5 (.A4( u1_u2_u2_n124 ) , .A3( u1_u2_u2_n125 ) , .A2( u1_u2_u2_n126 ) , .A1( u1_u2_u2_n127 ) , .ZN( u1_u2_u2_n128 ) );
  NAND2_X1 u1_u2_u2_U50 (.A1( u1_u2_u2_n100 ) , .A2( u1_u2_u2_n105 ) , .ZN( u1_u2_u2_n132 ) );
  INV_X1 u1_u2_u2_U51 (.A( u1_u2_u2_n140 ) , .ZN( u1_u2_u2_n168 ) );
  INV_X1 u1_u2_u2_U52 (.A( u1_u2_u2_n138 ) , .ZN( u1_u2_u2_n167 ) );
  OAI21_X1 u1_u2_u2_U53 (.A( u1_u2_u2_n141 ) , .B2( u1_u2_u2_n142 ) , .ZN( u1_u2_u2_n146 ) , .B1( u1_u2_u2_n153 ) );
  OAI21_X1 u1_u2_u2_U54 (.A( u1_u2_u2_n140 ) , .ZN( u1_u2_u2_n141 ) , .B1( u1_u2_u2_n176 ) , .B2( u1_u2_u2_n177 ) );
  NOR3_X1 u1_u2_u2_U55 (.ZN( u1_u2_u2_n142 ) , .A3( u1_u2_u2_n175 ) , .A2( u1_u2_u2_n178 ) , .A1( u1_u2_u2_n181 ) );
  NAND2_X1 u1_u2_u2_U56 (.A1( u1_u2_u2_n102 ) , .A2( u1_u2_u2_n106 ) , .ZN( u1_u2_u2_n113 ) );
  NAND2_X1 u1_u2_u2_U57 (.A1( u1_u2_u2_n106 ) , .A2( u1_u2_u2_n107 ) , .ZN( u1_u2_u2_n131 ) );
  NAND2_X1 u1_u2_u2_U58 (.A1( u1_u2_u2_n103 ) , .A2( u1_u2_u2_n107 ) , .ZN( u1_u2_u2_n139 ) );
  NAND2_X1 u1_u2_u2_U59 (.A1( u1_u2_u2_n103 ) , .A2( u1_u2_u2_n105 ) , .ZN( u1_u2_u2_n133 ) );
  AOI21_X1 u1_u2_u2_U6 (.B2( u1_u2_u2_n119 ) , .ZN( u1_u2_u2_n127 ) , .A( u1_u2_u2_n137 ) , .B1( u1_u2_u2_n155 ) );
  NAND2_X1 u1_u2_u2_U60 (.A1( u1_u2_u2_n102 ) , .A2( u1_u2_u2_n103 ) , .ZN( u1_u2_u2_n154 ) );
  NAND2_X1 u1_u2_u2_U61 (.A2( u1_u2_u2_n103 ) , .A1( u1_u2_u2_n104 ) , .ZN( u1_u2_u2_n119 ) );
  NAND2_X1 u1_u2_u2_U62 (.A2( u1_u2_u2_n107 ) , .A1( u1_u2_u2_n108 ) , .ZN( u1_u2_u2_n123 ) );
  NAND2_X1 u1_u2_u2_U63 (.A1( u1_u2_u2_n104 ) , .A2( u1_u2_u2_n108 ) , .ZN( u1_u2_u2_n122 ) );
  INV_X1 u1_u2_u2_U64 (.A( u1_u2_u2_n114 ) , .ZN( u1_u2_u2_n172 ) );
  NAND2_X1 u1_u2_u2_U65 (.A2( u1_u2_u2_n100 ) , .A1( u1_u2_u2_n102 ) , .ZN( u1_u2_u2_n116 ) );
  NAND2_X1 u1_u2_u2_U66 (.A1( u1_u2_u2_n102 ) , .A2( u1_u2_u2_n108 ) , .ZN( u1_u2_u2_n120 ) );
  NAND2_X1 u1_u2_u2_U67 (.A2( u1_u2_u2_n105 ) , .A1( u1_u2_u2_n106 ) , .ZN( u1_u2_u2_n117 ) );
  INV_X1 u1_u2_u2_U68 (.ZN( u1_u2_u2_n187 ) , .A( u1_u2_u2_n99 ) );
  OAI21_X1 u1_u2_u2_U69 (.B1( u1_u2_u2_n137 ) , .B2( u1_u2_u2_n143 ) , .A( u1_u2_u2_n98 ) , .ZN( u1_u2_u2_n99 ) );
  AOI21_X1 u1_u2_u2_U7 (.ZN( u1_u2_u2_n124 ) , .B1( u1_u2_u2_n131 ) , .B2( u1_u2_u2_n143 ) , .A( u1_u2_u2_n172 ) );
  NOR2_X1 u1_u2_u2_U70 (.A2( u1_u2_X_16 ) , .ZN( u1_u2_u2_n140 ) , .A1( u1_u2_u2_n166 ) );
  NOR2_X1 u1_u2_u2_U71 (.A2( u1_u2_X_13 ) , .A1( u1_u2_X_14 ) , .ZN( u1_u2_u2_n100 ) );
  NOR2_X1 u1_u2_u2_U72 (.A2( u1_u2_X_16 ) , .A1( u1_u2_X_17 ) , .ZN( u1_u2_u2_n138 ) );
  NOR2_X1 u1_u2_u2_U73 (.A2( u1_u2_X_15 ) , .A1( u1_u2_X_18 ) , .ZN( u1_u2_u2_n104 ) );
  NOR2_X1 u1_u2_u2_U74 (.A2( u1_u2_X_14 ) , .ZN( u1_u2_u2_n103 ) , .A1( u1_u2_u2_n174 ) );
  NOR2_X1 u1_u2_u2_U75 (.A2( u1_u2_X_15 ) , .ZN( u1_u2_u2_n102 ) , .A1( u1_u2_u2_n165 ) );
  NOR2_X1 u1_u2_u2_U76 (.A2( u1_u2_X_17 ) , .ZN( u1_u2_u2_n114 ) , .A1( u1_u2_u2_n169 ) );
  AND2_X1 u1_u2_u2_U77 (.A1( u1_u2_X_15 ) , .ZN( u1_u2_u2_n105 ) , .A2( u1_u2_u2_n165 ) );
  AND2_X1 u1_u2_u2_U78 (.A2( u1_u2_X_15 ) , .A1( u1_u2_X_18 ) , .ZN( u1_u2_u2_n107 ) );
  AND2_X1 u1_u2_u2_U79 (.A1( u1_u2_X_14 ) , .ZN( u1_u2_u2_n106 ) , .A2( u1_u2_u2_n174 ) );
  AOI21_X1 u1_u2_u2_U8 (.B2( u1_u2_u2_n120 ) , .B1( u1_u2_u2_n121 ) , .ZN( u1_u2_u2_n126 ) , .A( u1_u2_u2_n167 ) );
  AND2_X1 u1_u2_u2_U80 (.A1( u1_u2_X_13 ) , .A2( u1_u2_X_14 ) , .ZN( u1_u2_u2_n108 ) );
  INV_X1 u1_u2_u2_U81 (.A( u1_u2_X_16 ) , .ZN( u1_u2_u2_n169 ) );
  INV_X1 u1_u2_u2_U82 (.A( u1_u2_X_17 ) , .ZN( u1_u2_u2_n166 ) );
  INV_X1 u1_u2_u2_U83 (.A( u1_u2_X_13 ) , .ZN( u1_u2_u2_n174 ) );
  INV_X1 u1_u2_u2_U84 (.A( u1_u2_X_18 ) , .ZN( u1_u2_u2_n165 ) );
  NAND4_X1 u1_u2_u2_U85 (.ZN( u1_out2_24 ) , .A4( u1_u2_u2_n111 ) , .A3( u1_u2_u2_n112 ) , .A1( u1_u2_u2_n130 ) , .A2( u1_u2_u2_n187 ) );
  AOI21_X1 u1_u2_u2_U86 (.ZN( u1_u2_u2_n112 ) , .B2( u1_u2_u2_n156 ) , .A( u1_u2_u2_n164 ) , .B1( u1_u2_u2_n181 ) );
  AOI221_X1 u1_u2_u2_U87 (.A( u1_u2_u2_n109 ) , .B1( u1_u2_u2_n110 ) , .ZN( u1_u2_u2_n111 ) , .C1( u1_u2_u2_n134 ) , .C2( u1_u2_u2_n170 ) , .B2( u1_u2_u2_n173 ) );
  NAND4_X1 u1_u2_u2_U88 (.ZN( u1_out2_16 ) , .A4( u1_u2_u2_n128 ) , .A3( u1_u2_u2_n129 ) , .A1( u1_u2_u2_n130 ) , .A2( u1_u2_u2_n186 ) );
  AOI22_X1 u1_u2_u2_U89 (.A2( u1_u2_u2_n118 ) , .ZN( u1_u2_u2_n129 ) , .A1( u1_u2_u2_n140 ) , .B1( u1_u2_u2_n157 ) , .B2( u1_u2_u2_n170 ) );
  OAI22_X1 u1_u2_u2_U9 (.ZN( u1_u2_u2_n109 ) , .A2( u1_u2_u2_n113 ) , .B2( u1_u2_u2_n133 ) , .B1( u1_u2_u2_n167 ) , .A1( u1_u2_u2_n168 ) );
  INV_X1 u1_u2_u2_U90 (.A( u1_u2_u2_n163 ) , .ZN( u1_u2_u2_n186 ) );
  NAND4_X1 u1_u2_u2_U91 (.ZN( u1_out2_30 ) , .A4( u1_u2_u2_n147 ) , .A3( u1_u2_u2_n148 ) , .A2( u1_u2_u2_n149 ) , .A1( u1_u2_u2_n187 ) );
  NOR3_X1 u1_u2_u2_U92 (.A3( u1_u2_u2_n144 ) , .A2( u1_u2_u2_n145 ) , .A1( u1_u2_u2_n146 ) , .ZN( u1_u2_u2_n147 ) );
  AOI21_X1 u1_u2_u2_U93 (.B2( u1_u2_u2_n138 ) , .ZN( u1_u2_u2_n148 ) , .A( u1_u2_u2_n162 ) , .B1( u1_u2_u2_n182 ) );
  OR4_X1 u1_u2_u2_U94 (.ZN( u1_out2_6 ) , .A4( u1_u2_u2_n161 ) , .A3( u1_u2_u2_n162 ) , .A2( u1_u2_u2_n163 ) , .A1( u1_u2_u2_n164 ) );
  OR3_X1 u1_u2_u2_U95 (.A2( u1_u2_u2_n159 ) , .A1( u1_u2_u2_n160 ) , .ZN( u1_u2_u2_n161 ) , .A3( u1_u2_u2_n183 ) );
  AOI21_X1 u1_u2_u2_U96 (.B2( u1_u2_u2_n154 ) , .B1( u1_u2_u2_n155 ) , .ZN( u1_u2_u2_n159 ) , .A( u1_u2_u2_n167 ) );
  NAND3_X1 u1_u2_u2_U97 (.A2( u1_u2_u2_n117 ) , .A1( u1_u2_u2_n122 ) , .A3( u1_u2_u2_n123 ) , .ZN( u1_u2_u2_n134 ) );
  NAND3_X1 u1_u2_u2_U98 (.ZN( u1_u2_u2_n110 ) , .A2( u1_u2_u2_n131 ) , .A3( u1_u2_u2_n139 ) , .A1( u1_u2_u2_n154 ) );
  NAND3_X1 u1_u2_u2_U99 (.A2( u1_u2_u2_n100 ) , .ZN( u1_u2_u2_n101 ) , .A1( u1_u2_u2_n104 ) , .A3( u1_u2_u2_n114 ) );
  OAI22_X1 u1_u2_u3_U10 (.B1( u1_u2_u3_n113 ) , .A2( u1_u2_u3_n135 ) , .A1( u1_u2_u3_n150 ) , .B2( u1_u2_u3_n164 ) , .ZN( u1_u2_u3_n98 ) );
  OAI211_X1 u1_u2_u3_U11 (.B( u1_u2_u3_n106 ) , .ZN( u1_u2_u3_n119 ) , .C2( u1_u2_u3_n128 ) , .C1( u1_u2_u3_n167 ) , .A( u1_u2_u3_n181 ) );
  AOI221_X1 u1_u2_u3_U12 (.C1( u1_u2_u3_n105 ) , .ZN( u1_u2_u3_n106 ) , .A( u1_u2_u3_n131 ) , .B2( u1_u2_u3_n132 ) , .C2( u1_u2_u3_n133 ) , .B1( u1_u2_u3_n169 ) );
  INV_X1 u1_u2_u3_U13 (.ZN( u1_u2_u3_n181 ) , .A( u1_u2_u3_n98 ) );
  NAND2_X1 u1_u2_u3_U14 (.ZN( u1_u2_u3_n105 ) , .A2( u1_u2_u3_n130 ) , .A1( u1_u2_u3_n155 ) );
  AOI22_X1 u1_u2_u3_U15 (.B1( u1_u2_u3_n115 ) , .A2( u1_u2_u3_n116 ) , .ZN( u1_u2_u3_n123 ) , .B2( u1_u2_u3_n133 ) , .A1( u1_u2_u3_n169 ) );
  NAND2_X1 u1_u2_u3_U16 (.ZN( u1_u2_u3_n116 ) , .A2( u1_u2_u3_n151 ) , .A1( u1_u2_u3_n182 ) );
  NOR2_X1 u1_u2_u3_U17 (.ZN( u1_u2_u3_n126 ) , .A2( u1_u2_u3_n150 ) , .A1( u1_u2_u3_n164 ) );
  AOI21_X1 u1_u2_u3_U18 (.ZN( u1_u2_u3_n112 ) , .B2( u1_u2_u3_n146 ) , .B1( u1_u2_u3_n155 ) , .A( u1_u2_u3_n167 ) );
  NAND2_X1 u1_u2_u3_U19 (.A1( u1_u2_u3_n135 ) , .ZN( u1_u2_u3_n142 ) , .A2( u1_u2_u3_n164 ) );
  NAND2_X1 u1_u2_u3_U20 (.ZN( u1_u2_u3_n132 ) , .A2( u1_u2_u3_n152 ) , .A1( u1_u2_u3_n156 ) );
  AND2_X1 u1_u2_u3_U21 (.A2( u1_u2_u3_n113 ) , .A1( u1_u2_u3_n114 ) , .ZN( u1_u2_u3_n151 ) );
  INV_X1 u1_u2_u3_U22 (.A( u1_u2_u3_n133 ) , .ZN( u1_u2_u3_n165 ) );
  INV_X1 u1_u2_u3_U23 (.A( u1_u2_u3_n135 ) , .ZN( u1_u2_u3_n170 ) );
  NAND2_X1 u1_u2_u3_U24 (.A1( u1_u2_u3_n107 ) , .A2( u1_u2_u3_n108 ) , .ZN( u1_u2_u3_n140 ) );
  NAND2_X1 u1_u2_u3_U25 (.ZN( u1_u2_u3_n117 ) , .A1( u1_u2_u3_n124 ) , .A2( u1_u2_u3_n148 ) );
  NAND2_X1 u1_u2_u3_U26 (.ZN( u1_u2_u3_n143 ) , .A1( u1_u2_u3_n165 ) , .A2( u1_u2_u3_n167 ) );
  INV_X1 u1_u2_u3_U27 (.A( u1_u2_u3_n130 ) , .ZN( u1_u2_u3_n177 ) );
  INV_X1 u1_u2_u3_U28 (.A( u1_u2_u3_n128 ) , .ZN( u1_u2_u3_n176 ) );
  INV_X1 u1_u2_u3_U29 (.A( u1_u2_u3_n155 ) , .ZN( u1_u2_u3_n174 ) );
  INV_X1 u1_u2_u3_U3 (.A( u1_u2_u3_n129 ) , .ZN( u1_u2_u3_n183 ) );
  INV_X1 u1_u2_u3_U30 (.A( u1_u2_u3_n139 ) , .ZN( u1_u2_u3_n185 ) );
  NOR2_X1 u1_u2_u3_U31 (.ZN( u1_u2_u3_n135 ) , .A2( u1_u2_u3_n141 ) , .A1( u1_u2_u3_n169 ) );
  OAI222_X1 u1_u2_u3_U32 (.C2( u1_u2_u3_n107 ) , .A2( u1_u2_u3_n108 ) , .B1( u1_u2_u3_n135 ) , .ZN( u1_u2_u3_n138 ) , .B2( u1_u2_u3_n146 ) , .C1( u1_u2_u3_n154 ) , .A1( u1_u2_u3_n164 ) );
  NOR4_X1 u1_u2_u3_U33 (.A4( u1_u2_u3_n157 ) , .A3( u1_u2_u3_n158 ) , .A2( u1_u2_u3_n159 ) , .A1( u1_u2_u3_n160 ) , .ZN( u1_u2_u3_n161 ) );
  AOI21_X1 u1_u2_u3_U34 (.B2( u1_u2_u3_n152 ) , .B1( u1_u2_u3_n153 ) , .ZN( u1_u2_u3_n158 ) , .A( u1_u2_u3_n164 ) );
  AOI21_X1 u1_u2_u3_U35 (.A( u1_u2_u3_n154 ) , .B2( u1_u2_u3_n155 ) , .B1( u1_u2_u3_n156 ) , .ZN( u1_u2_u3_n157 ) );
  AOI21_X1 u1_u2_u3_U36 (.A( u1_u2_u3_n149 ) , .B2( u1_u2_u3_n150 ) , .B1( u1_u2_u3_n151 ) , .ZN( u1_u2_u3_n159 ) );
  AOI211_X1 u1_u2_u3_U37 (.ZN( u1_u2_u3_n109 ) , .A( u1_u2_u3_n119 ) , .C2( u1_u2_u3_n129 ) , .B( u1_u2_u3_n138 ) , .C1( u1_u2_u3_n141 ) );
  AOI211_X1 u1_u2_u3_U38 (.B( u1_u2_u3_n119 ) , .A( u1_u2_u3_n120 ) , .C2( u1_u2_u3_n121 ) , .ZN( u1_u2_u3_n122 ) , .C1( u1_u2_u3_n179 ) );
  INV_X1 u1_u2_u3_U39 (.A( u1_u2_u3_n156 ) , .ZN( u1_u2_u3_n179 ) );
  INV_X1 u1_u2_u3_U4 (.A( u1_u2_u3_n140 ) , .ZN( u1_u2_u3_n182 ) );
  OAI22_X1 u1_u2_u3_U40 (.B1( u1_u2_u3_n118 ) , .ZN( u1_u2_u3_n120 ) , .A1( u1_u2_u3_n135 ) , .B2( u1_u2_u3_n154 ) , .A2( u1_u2_u3_n178 ) );
  AND3_X1 u1_u2_u3_U41 (.ZN( u1_u2_u3_n118 ) , .A2( u1_u2_u3_n124 ) , .A1( u1_u2_u3_n144 ) , .A3( u1_u2_u3_n152 ) );
  INV_X1 u1_u2_u3_U42 (.A( u1_u2_u3_n121 ) , .ZN( u1_u2_u3_n164 ) );
  NAND2_X1 u1_u2_u3_U43 (.ZN( u1_u2_u3_n133 ) , .A1( u1_u2_u3_n154 ) , .A2( u1_u2_u3_n164 ) );
  OAI211_X1 u1_u2_u3_U44 (.B( u1_u2_u3_n127 ) , .ZN( u1_u2_u3_n139 ) , .C1( u1_u2_u3_n150 ) , .C2( u1_u2_u3_n154 ) , .A( u1_u2_u3_n184 ) );
  INV_X1 u1_u2_u3_U45 (.A( u1_u2_u3_n125 ) , .ZN( u1_u2_u3_n184 ) );
  AOI221_X1 u1_u2_u3_U46 (.A( u1_u2_u3_n126 ) , .ZN( u1_u2_u3_n127 ) , .C2( u1_u2_u3_n132 ) , .C1( u1_u2_u3_n169 ) , .B2( u1_u2_u3_n170 ) , .B1( u1_u2_u3_n174 ) );
  OAI22_X1 u1_u2_u3_U47 (.A1( u1_u2_u3_n124 ) , .ZN( u1_u2_u3_n125 ) , .B2( u1_u2_u3_n145 ) , .A2( u1_u2_u3_n165 ) , .B1( u1_u2_u3_n167 ) );
  NOR2_X1 u1_u2_u3_U48 (.A1( u1_u2_u3_n113 ) , .ZN( u1_u2_u3_n131 ) , .A2( u1_u2_u3_n154 ) );
  NAND2_X1 u1_u2_u3_U49 (.A1( u1_u2_u3_n103 ) , .ZN( u1_u2_u3_n150 ) , .A2( u1_u2_u3_n99 ) );
  INV_X1 u1_u2_u3_U5 (.A( u1_u2_u3_n117 ) , .ZN( u1_u2_u3_n178 ) );
  NAND2_X1 u1_u2_u3_U50 (.A2( u1_u2_u3_n102 ) , .ZN( u1_u2_u3_n155 ) , .A1( u1_u2_u3_n97 ) );
  INV_X1 u1_u2_u3_U51 (.A( u1_u2_u3_n141 ) , .ZN( u1_u2_u3_n167 ) );
  AOI21_X1 u1_u2_u3_U52 (.B2( u1_u2_u3_n114 ) , .B1( u1_u2_u3_n146 ) , .A( u1_u2_u3_n154 ) , .ZN( u1_u2_u3_n94 ) );
  AOI21_X1 u1_u2_u3_U53 (.ZN( u1_u2_u3_n110 ) , .B2( u1_u2_u3_n142 ) , .B1( u1_u2_u3_n186 ) , .A( u1_u2_u3_n95 ) );
  INV_X1 u1_u2_u3_U54 (.A( u1_u2_u3_n145 ) , .ZN( u1_u2_u3_n186 ) );
  AOI21_X1 u1_u2_u3_U55 (.B1( u1_u2_u3_n124 ) , .A( u1_u2_u3_n149 ) , .B2( u1_u2_u3_n155 ) , .ZN( u1_u2_u3_n95 ) );
  INV_X1 u1_u2_u3_U56 (.A( u1_u2_u3_n149 ) , .ZN( u1_u2_u3_n169 ) );
  NAND2_X1 u1_u2_u3_U57 (.ZN( u1_u2_u3_n124 ) , .A1( u1_u2_u3_n96 ) , .A2( u1_u2_u3_n97 ) );
  NAND2_X1 u1_u2_u3_U58 (.A2( u1_u2_u3_n100 ) , .ZN( u1_u2_u3_n146 ) , .A1( u1_u2_u3_n96 ) );
  NAND2_X1 u1_u2_u3_U59 (.A1( u1_u2_u3_n101 ) , .ZN( u1_u2_u3_n145 ) , .A2( u1_u2_u3_n99 ) );
  AOI221_X1 u1_u2_u3_U6 (.A( u1_u2_u3_n131 ) , .C2( u1_u2_u3_n132 ) , .C1( u1_u2_u3_n133 ) , .ZN( u1_u2_u3_n134 ) , .B1( u1_u2_u3_n143 ) , .B2( u1_u2_u3_n177 ) );
  NAND2_X1 u1_u2_u3_U60 (.A1( u1_u2_u3_n100 ) , .ZN( u1_u2_u3_n156 ) , .A2( u1_u2_u3_n99 ) );
  NAND2_X1 u1_u2_u3_U61 (.A2( u1_u2_u3_n101 ) , .A1( u1_u2_u3_n104 ) , .ZN( u1_u2_u3_n148 ) );
  NAND2_X1 u1_u2_u3_U62 (.A1( u1_u2_u3_n100 ) , .A2( u1_u2_u3_n102 ) , .ZN( u1_u2_u3_n128 ) );
  NAND2_X1 u1_u2_u3_U63 (.A2( u1_u2_u3_n101 ) , .A1( u1_u2_u3_n102 ) , .ZN( u1_u2_u3_n152 ) );
  NAND2_X1 u1_u2_u3_U64 (.A2( u1_u2_u3_n101 ) , .ZN( u1_u2_u3_n114 ) , .A1( u1_u2_u3_n96 ) );
  NAND2_X1 u1_u2_u3_U65 (.ZN( u1_u2_u3_n107 ) , .A1( u1_u2_u3_n97 ) , .A2( u1_u2_u3_n99 ) );
  NAND2_X1 u1_u2_u3_U66 (.A2( u1_u2_u3_n100 ) , .A1( u1_u2_u3_n104 ) , .ZN( u1_u2_u3_n113 ) );
  NAND2_X1 u1_u2_u3_U67 (.A1( u1_u2_u3_n104 ) , .ZN( u1_u2_u3_n153 ) , .A2( u1_u2_u3_n97 ) );
  NAND2_X1 u1_u2_u3_U68 (.A2( u1_u2_u3_n103 ) , .A1( u1_u2_u3_n104 ) , .ZN( u1_u2_u3_n130 ) );
  NAND2_X1 u1_u2_u3_U69 (.A2( u1_u2_u3_n103 ) , .ZN( u1_u2_u3_n144 ) , .A1( u1_u2_u3_n96 ) );
  OAI22_X1 u1_u2_u3_U7 (.B2( u1_u2_u3_n147 ) , .A2( u1_u2_u3_n148 ) , .ZN( u1_u2_u3_n160 ) , .B1( u1_u2_u3_n165 ) , .A1( u1_u2_u3_n168 ) );
  NAND2_X1 u1_u2_u3_U70 (.A1( u1_u2_u3_n102 ) , .A2( u1_u2_u3_n103 ) , .ZN( u1_u2_u3_n108 ) );
  NOR2_X1 u1_u2_u3_U71 (.A2( u1_u2_X_19 ) , .A1( u1_u2_X_20 ) , .ZN( u1_u2_u3_n99 ) );
  NOR2_X1 u1_u2_u3_U72 (.A2( u1_u2_X_21 ) , .A1( u1_u2_X_24 ) , .ZN( u1_u2_u3_n103 ) );
  NOR2_X1 u1_u2_u3_U73 (.A2( u1_u2_X_24 ) , .A1( u1_u2_u3_n171 ) , .ZN( u1_u2_u3_n97 ) );
  NOR2_X1 u1_u2_u3_U74 (.A2( u1_u2_X_23 ) , .ZN( u1_u2_u3_n141 ) , .A1( u1_u2_u3_n166 ) );
  NOR2_X1 u1_u2_u3_U75 (.A2( u1_u2_X_19 ) , .A1( u1_u2_u3_n172 ) , .ZN( u1_u2_u3_n96 ) );
  NAND2_X1 u1_u2_u3_U76 (.A1( u1_u2_X_22 ) , .A2( u1_u2_X_23 ) , .ZN( u1_u2_u3_n154 ) );
  NAND2_X1 u1_u2_u3_U77 (.A1( u1_u2_X_23 ) , .ZN( u1_u2_u3_n149 ) , .A2( u1_u2_u3_n166 ) );
  NOR2_X1 u1_u2_u3_U78 (.A2( u1_u2_X_22 ) , .A1( u1_u2_X_23 ) , .ZN( u1_u2_u3_n121 ) );
  AND2_X1 u1_u2_u3_U79 (.A1( u1_u2_X_24 ) , .ZN( u1_u2_u3_n101 ) , .A2( u1_u2_u3_n171 ) );
  AND3_X1 u1_u2_u3_U8 (.A3( u1_u2_u3_n144 ) , .A2( u1_u2_u3_n145 ) , .A1( u1_u2_u3_n146 ) , .ZN( u1_u2_u3_n147 ) );
  AND2_X1 u1_u2_u3_U80 (.A1( u1_u2_X_19 ) , .ZN( u1_u2_u3_n102 ) , .A2( u1_u2_u3_n172 ) );
  AND2_X1 u1_u2_u3_U81 (.A1( u1_u2_X_21 ) , .A2( u1_u2_X_24 ) , .ZN( u1_u2_u3_n100 ) );
  AND2_X1 u1_u2_u3_U82 (.A2( u1_u2_X_19 ) , .A1( u1_u2_X_20 ) , .ZN( u1_u2_u3_n104 ) );
  INV_X1 u1_u2_u3_U83 (.A( u1_u2_X_22 ) , .ZN( u1_u2_u3_n166 ) );
  INV_X1 u1_u2_u3_U84 (.A( u1_u2_X_21 ) , .ZN( u1_u2_u3_n171 ) );
  INV_X1 u1_u2_u3_U85 (.A( u1_u2_X_20 ) , .ZN( u1_u2_u3_n172 ) );
  OR4_X1 u1_u2_u3_U86 (.ZN( u1_out2_10 ) , .A4( u1_u2_u3_n136 ) , .A3( u1_u2_u3_n137 ) , .A1( u1_u2_u3_n138 ) , .A2( u1_u2_u3_n139 ) );
  OAI222_X1 u1_u2_u3_U87 (.C1( u1_u2_u3_n128 ) , .ZN( u1_u2_u3_n137 ) , .B1( u1_u2_u3_n148 ) , .A2( u1_u2_u3_n150 ) , .B2( u1_u2_u3_n154 ) , .C2( u1_u2_u3_n164 ) , .A1( u1_u2_u3_n167 ) );
  OAI221_X1 u1_u2_u3_U88 (.A( u1_u2_u3_n134 ) , .B2( u1_u2_u3_n135 ) , .ZN( u1_u2_u3_n136 ) , .C1( u1_u2_u3_n149 ) , .B1( u1_u2_u3_n151 ) , .C2( u1_u2_u3_n183 ) );
  NAND4_X1 u1_u2_u3_U89 (.ZN( u1_out2_26 ) , .A4( u1_u2_u3_n109 ) , .A3( u1_u2_u3_n110 ) , .A2( u1_u2_u3_n111 ) , .A1( u1_u2_u3_n173 ) );
  INV_X1 u1_u2_u3_U9 (.A( u1_u2_u3_n143 ) , .ZN( u1_u2_u3_n168 ) );
  INV_X1 u1_u2_u3_U90 (.ZN( u1_u2_u3_n173 ) , .A( u1_u2_u3_n94 ) );
  OAI21_X1 u1_u2_u3_U91 (.ZN( u1_u2_u3_n111 ) , .B2( u1_u2_u3_n117 ) , .A( u1_u2_u3_n133 ) , .B1( u1_u2_u3_n176 ) );
  NAND4_X1 u1_u2_u3_U92 (.ZN( u1_out2_20 ) , .A4( u1_u2_u3_n122 ) , .A3( u1_u2_u3_n123 ) , .A1( u1_u2_u3_n175 ) , .A2( u1_u2_u3_n180 ) );
  INV_X1 u1_u2_u3_U93 (.A( u1_u2_u3_n112 ) , .ZN( u1_u2_u3_n175 ) );
  INV_X1 u1_u2_u3_U94 (.A( u1_u2_u3_n126 ) , .ZN( u1_u2_u3_n180 ) );
  NAND4_X1 u1_u2_u3_U95 (.ZN( u1_out2_1 ) , .A4( u1_u2_u3_n161 ) , .A3( u1_u2_u3_n162 ) , .A2( u1_u2_u3_n163 ) , .A1( u1_u2_u3_n185 ) );
  NAND2_X1 u1_u2_u3_U96 (.ZN( u1_u2_u3_n163 ) , .A2( u1_u2_u3_n170 ) , .A1( u1_u2_u3_n176 ) );
  AOI22_X1 u1_u2_u3_U97 (.B2( u1_u2_u3_n140 ) , .B1( u1_u2_u3_n141 ) , .A2( u1_u2_u3_n142 ) , .ZN( u1_u2_u3_n162 ) , .A1( u1_u2_u3_n177 ) );
  NAND3_X1 u1_u2_u3_U98 (.A1( u1_u2_u3_n114 ) , .ZN( u1_u2_u3_n115 ) , .A2( u1_u2_u3_n145 ) , .A3( u1_u2_u3_n153 ) );
  NAND3_X1 u1_u2_u3_U99 (.ZN( u1_u2_u3_n129 ) , .A2( u1_u2_u3_n144 ) , .A1( u1_u2_u3_n153 ) , .A3( u1_u2_u3_n182 ) );
  XOR2_X1 u1_u4_U16 (.B( u1_K5_3 ) , .A( u1_R3_2 ) , .Z( u1_u4_X_3 ) );
  XOR2_X1 u1_u4_U27 (.B( u1_K5_2 ) , .A( u1_R3_1 ) , .Z( u1_u4_X_2 ) );
  XOR2_X1 u1_u4_U38 (.B( u1_K5_1 ) , .A( u1_R3_32 ) , .Z( u1_u4_X_1 ) );
  XOR2_X1 u1_u4_U4 (.B( u1_K5_6 ) , .A( u1_R3_5 ) , .Z( u1_u4_X_6 ) );
  XOR2_X1 u1_u4_U40 (.B( u1_K5_18 ) , .A( u1_R3_13 ) , .Z( u1_u4_X_18 ) );
  XOR2_X1 u1_u4_U41 (.B( u1_K5_17 ) , .A( u1_R3_12 ) , .Z( u1_u4_X_17 ) );
  XOR2_X1 u1_u4_U42 (.B( u1_K5_16 ) , .A( u1_R3_11 ) , .Z( u1_u4_X_16 ) );
  XOR2_X1 u1_u4_U43 (.B( u1_K5_15 ) , .A( u1_R3_10 ) , .Z( u1_u4_X_15 ) );
  XOR2_X1 u1_u4_U44 (.B( u1_K5_14 ) , .A( u1_R3_9 ) , .Z( u1_u4_X_14 ) );
  XOR2_X1 u1_u4_U45 (.B( u1_K5_13 ) , .A( u1_R3_8 ) , .Z( u1_u4_X_13 ) );
  XOR2_X1 u1_u4_U5 (.B( u1_K5_5 ) , .A( u1_R3_4 ) , .Z( u1_u4_X_5 ) );
  XOR2_X1 u1_u4_U6 (.B( u1_K5_4 ) , .A( u1_R3_3 ) , .Z( u1_u4_X_4 ) );
  AND3_X1 u1_u4_u0_U10 (.A2( u1_u4_u0_n112 ) , .ZN( u1_u4_u0_n127 ) , .A3( u1_u4_u0_n130 ) , .A1( u1_u4_u0_n148 ) );
  NAND2_X1 u1_u4_u0_U11 (.ZN( u1_u4_u0_n113 ) , .A1( u1_u4_u0_n139 ) , .A2( u1_u4_u0_n149 ) );
  AND2_X1 u1_u4_u0_U12 (.ZN( u1_u4_u0_n107 ) , .A1( u1_u4_u0_n130 ) , .A2( u1_u4_u0_n140 ) );
  AND2_X1 u1_u4_u0_U13 (.A2( u1_u4_u0_n129 ) , .A1( u1_u4_u0_n130 ) , .ZN( u1_u4_u0_n151 ) );
  AND2_X1 u1_u4_u0_U14 (.A1( u1_u4_u0_n108 ) , .A2( u1_u4_u0_n125 ) , .ZN( u1_u4_u0_n145 ) );
  INV_X1 u1_u4_u0_U15 (.A( u1_u4_u0_n143 ) , .ZN( u1_u4_u0_n173 ) );
  NOR2_X1 u1_u4_u0_U16 (.A2( u1_u4_u0_n136 ) , .ZN( u1_u4_u0_n147 ) , .A1( u1_u4_u0_n160 ) );
  NOR2_X1 u1_u4_u0_U17 (.A1( u1_u4_u0_n163 ) , .A2( u1_u4_u0_n164 ) , .ZN( u1_u4_u0_n95 ) );
  AOI21_X1 u1_u4_u0_U18 (.B1( u1_u4_u0_n103 ) , .ZN( u1_u4_u0_n132 ) , .A( u1_u4_u0_n165 ) , .B2( u1_u4_u0_n93 ) );
  INV_X1 u1_u4_u0_U19 (.A( u1_u4_u0_n142 ) , .ZN( u1_u4_u0_n165 ) );
  OAI221_X1 u1_u4_u0_U20 (.C1( u1_u4_u0_n112 ) , .ZN( u1_u4_u0_n120 ) , .B1( u1_u4_u0_n138 ) , .B2( u1_u4_u0_n141 ) , .C2( u1_u4_u0_n147 ) , .A( u1_u4_u0_n172 ) );
  AOI211_X1 u1_u4_u0_U21 (.B( u1_u4_u0_n115 ) , .A( u1_u4_u0_n116 ) , .C2( u1_u4_u0_n117 ) , .C1( u1_u4_u0_n118 ) , .ZN( u1_u4_u0_n119 ) );
  OAI22_X1 u1_u4_u0_U22 (.B1( u1_u4_u0_n125 ) , .ZN( u1_u4_u0_n126 ) , .A1( u1_u4_u0_n138 ) , .A2( u1_u4_u0_n146 ) , .B2( u1_u4_u0_n147 ) );
  OAI22_X1 u1_u4_u0_U23 (.B1( u1_u4_u0_n131 ) , .A1( u1_u4_u0_n144 ) , .B2( u1_u4_u0_n147 ) , .A2( u1_u4_u0_n90 ) , .ZN( u1_u4_u0_n91 ) );
  AND3_X1 u1_u4_u0_U24 (.A3( u1_u4_u0_n121 ) , .A2( u1_u4_u0_n125 ) , .A1( u1_u4_u0_n148 ) , .ZN( u1_u4_u0_n90 ) );
  INV_X1 u1_u4_u0_U25 (.A( u1_u4_u0_n136 ) , .ZN( u1_u4_u0_n161 ) );
  AOI22_X1 u1_u4_u0_U26 (.B2( u1_u4_u0_n109 ) , .A2( u1_u4_u0_n110 ) , .ZN( u1_u4_u0_n111 ) , .B1( u1_u4_u0_n118 ) , .A1( u1_u4_u0_n160 ) );
  INV_X1 u1_u4_u0_U27 (.A( u1_u4_u0_n118 ) , .ZN( u1_u4_u0_n158 ) );
  AOI21_X1 u1_u4_u0_U28 (.ZN( u1_u4_u0_n104 ) , .B1( u1_u4_u0_n107 ) , .B2( u1_u4_u0_n141 ) , .A( u1_u4_u0_n144 ) );
  AOI21_X1 u1_u4_u0_U29 (.B1( u1_u4_u0_n127 ) , .B2( u1_u4_u0_n129 ) , .A( u1_u4_u0_n138 ) , .ZN( u1_u4_u0_n96 ) );
  INV_X1 u1_u4_u0_U3 (.A( u1_u4_u0_n113 ) , .ZN( u1_u4_u0_n166 ) );
  AOI21_X1 u1_u4_u0_U30 (.ZN( u1_u4_u0_n116 ) , .B2( u1_u4_u0_n142 ) , .A( u1_u4_u0_n144 ) , .B1( u1_u4_u0_n166 ) );
  NAND2_X1 u1_u4_u0_U31 (.A1( u1_u4_u0_n100 ) , .A2( u1_u4_u0_n103 ) , .ZN( u1_u4_u0_n125 ) );
  NAND2_X1 u1_u4_u0_U32 (.A1( u1_u4_u0_n101 ) , .A2( u1_u4_u0_n102 ) , .ZN( u1_u4_u0_n150 ) );
  INV_X1 u1_u4_u0_U33 (.A( u1_u4_u0_n138 ) , .ZN( u1_u4_u0_n160 ) );
  NAND2_X1 u1_u4_u0_U34 (.A1( u1_u4_u0_n102 ) , .ZN( u1_u4_u0_n128 ) , .A2( u1_u4_u0_n95 ) );
  NAND2_X1 u1_u4_u0_U35 (.A1( u1_u4_u0_n100 ) , .ZN( u1_u4_u0_n129 ) , .A2( u1_u4_u0_n95 ) );
  NAND2_X1 u1_u4_u0_U36 (.A2( u1_u4_u0_n100 ) , .ZN( u1_u4_u0_n131 ) , .A1( u1_u4_u0_n92 ) );
  NAND2_X1 u1_u4_u0_U37 (.A2( u1_u4_u0_n100 ) , .A1( u1_u4_u0_n101 ) , .ZN( u1_u4_u0_n139 ) );
  NAND2_X1 u1_u4_u0_U38 (.ZN( u1_u4_u0_n148 ) , .A1( u1_u4_u0_n93 ) , .A2( u1_u4_u0_n95 ) );
  NAND2_X1 u1_u4_u0_U39 (.A2( u1_u4_u0_n102 ) , .A1( u1_u4_u0_n103 ) , .ZN( u1_u4_u0_n149 ) );
  AOI21_X1 u1_u4_u0_U4 (.B1( u1_u4_u0_n114 ) , .ZN( u1_u4_u0_n115 ) , .B2( u1_u4_u0_n129 ) , .A( u1_u4_u0_n161 ) );
  NAND2_X1 u1_u4_u0_U40 (.A2( u1_u4_u0_n102 ) , .ZN( u1_u4_u0_n114 ) , .A1( u1_u4_u0_n92 ) );
  NAND2_X1 u1_u4_u0_U41 (.A2( u1_u4_u0_n101 ) , .ZN( u1_u4_u0_n121 ) , .A1( u1_u4_u0_n93 ) );
  INV_X1 u1_u4_u0_U42 (.ZN( u1_u4_u0_n172 ) , .A( u1_u4_u0_n88 ) );
  OAI222_X1 u1_u4_u0_U43 (.C1( u1_u4_u0_n108 ) , .A1( u1_u4_u0_n125 ) , .B2( u1_u4_u0_n128 ) , .B1( u1_u4_u0_n144 ) , .A2( u1_u4_u0_n158 ) , .C2( u1_u4_u0_n161 ) , .ZN( u1_u4_u0_n88 ) );
  NAND2_X1 u1_u4_u0_U44 (.ZN( u1_u4_u0_n112 ) , .A2( u1_u4_u0_n92 ) , .A1( u1_u4_u0_n93 ) );
  OR3_X1 u1_u4_u0_U45 (.A3( u1_u4_u0_n152 ) , .A2( u1_u4_u0_n153 ) , .A1( u1_u4_u0_n154 ) , .ZN( u1_u4_u0_n155 ) );
  AOI21_X1 u1_u4_u0_U46 (.A( u1_u4_u0_n144 ) , .B2( u1_u4_u0_n145 ) , .B1( u1_u4_u0_n146 ) , .ZN( u1_u4_u0_n154 ) );
  AOI21_X1 u1_u4_u0_U47 (.B2( u1_u4_u0_n150 ) , .B1( u1_u4_u0_n151 ) , .ZN( u1_u4_u0_n152 ) , .A( u1_u4_u0_n158 ) );
  AOI21_X1 u1_u4_u0_U48 (.A( u1_u4_u0_n147 ) , .B2( u1_u4_u0_n148 ) , .B1( u1_u4_u0_n149 ) , .ZN( u1_u4_u0_n153 ) );
  INV_X1 u1_u4_u0_U49 (.ZN( u1_u4_u0_n171 ) , .A( u1_u4_u0_n99 ) );
  AOI21_X1 u1_u4_u0_U5 (.B2( u1_u4_u0_n131 ) , .ZN( u1_u4_u0_n134 ) , .B1( u1_u4_u0_n151 ) , .A( u1_u4_u0_n158 ) );
  OAI211_X1 u1_u4_u0_U50 (.C2( u1_u4_u0_n140 ) , .C1( u1_u4_u0_n161 ) , .A( u1_u4_u0_n169 ) , .B( u1_u4_u0_n98 ) , .ZN( u1_u4_u0_n99 ) );
  INV_X1 u1_u4_u0_U51 (.ZN( u1_u4_u0_n169 ) , .A( u1_u4_u0_n91 ) );
  AOI211_X1 u1_u4_u0_U52 (.C1( u1_u4_u0_n118 ) , .A( u1_u4_u0_n123 ) , .B( u1_u4_u0_n96 ) , .C2( u1_u4_u0_n97 ) , .ZN( u1_u4_u0_n98 ) );
  NOR2_X1 u1_u4_u0_U53 (.A2( u1_u4_X_6 ) , .ZN( u1_u4_u0_n100 ) , .A1( u1_u4_u0_n162 ) );
  NOR2_X1 u1_u4_u0_U54 (.A2( u1_u4_X_4 ) , .A1( u1_u4_X_5 ) , .ZN( u1_u4_u0_n118 ) );
  NOR2_X1 u1_u4_u0_U55 (.A2( u1_u4_X_2 ) , .ZN( u1_u4_u0_n103 ) , .A1( u1_u4_u0_n164 ) );
  NOR2_X1 u1_u4_u0_U56 (.A2( u1_u4_X_1 ) , .A1( u1_u4_X_2 ) , .ZN( u1_u4_u0_n92 ) );
  NOR2_X1 u1_u4_u0_U57 (.A2( u1_u4_X_1 ) , .ZN( u1_u4_u0_n101 ) , .A1( u1_u4_u0_n163 ) );
  NAND2_X1 u1_u4_u0_U58 (.A2( u1_u4_X_4 ) , .A1( u1_u4_X_5 ) , .ZN( u1_u4_u0_n144 ) );
  NOR2_X1 u1_u4_u0_U59 (.A2( u1_u4_X_5 ) , .ZN( u1_u4_u0_n136 ) , .A1( u1_u4_u0_n159 ) );
  NOR2_X1 u1_u4_u0_U6 (.A1( u1_u4_u0_n108 ) , .ZN( u1_u4_u0_n123 ) , .A2( u1_u4_u0_n158 ) );
  NAND2_X1 u1_u4_u0_U60 (.A1( u1_u4_X_5 ) , .ZN( u1_u4_u0_n138 ) , .A2( u1_u4_u0_n159 ) );
  NOR2_X1 u1_u4_u0_U61 (.A2( u1_u4_X_3 ) , .A1( u1_u4_X_6 ) , .ZN( u1_u4_u0_n94 ) );
  AND2_X1 u1_u4_u0_U62 (.A2( u1_u4_X_3 ) , .A1( u1_u4_X_6 ) , .ZN( u1_u4_u0_n102 ) );
  AND2_X1 u1_u4_u0_U63 (.A1( u1_u4_X_6 ) , .A2( u1_u4_u0_n162 ) , .ZN( u1_u4_u0_n93 ) );
  INV_X1 u1_u4_u0_U64 (.A( u1_u4_X_4 ) , .ZN( u1_u4_u0_n159 ) );
  INV_X1 u1_u4_u0_U65 (.A( u1_u4_X_1 ) , .ZN( u1_u4_u0_n164 ) );
  INV_X1 u1_u4_u0_U66 (.A( u1_u4_X_2 ) , .ZN( u1_u4_u0_n163 ) );
  INV_X1 u1_u4_u0_U67 (.A( u1_u4_X_3 ) , .ZN( u1_u4_u0_n162 ) );
  INV_X1 u1_u4_u0_U68 (.A( u1_u4_u0_n126 ) , .ZN( u1_u4_u0_n168 ) );
  AOI211_X1 u1_u4_u0_U69 (.B( u1_u4_u0_n133 ) , .A( u1_u4_u0_n134 ) , .C2( u1_u4_u0_n135 ) , .C1( u1_u4_u0_n136 ) , .ZN( u1_u4_u0_n137 ) );
  OAI21_X1 u1_u4_u0_U7 (.B1( u1_u4_u0_n150 ) , .B2( u1_u4_u0_n158 ) , .A( u1_u4_u0_n172 ) , .ZN( u1_u4_u0_n89 ) );
  AOI21_X1 u1_u4_u0_U70 (.B2( u1_u4_u0_n107 ) , .ZN( u1_u4_u0_n124 ) , .B1( u1_u4_u0_n128 ) , .A( u1_u4_u0_n161 ) );
  INV_X1 u1_u4_u0_U71 (.A( u1_u4_u0_n111 ) , .ZN( u1_u4_u0_n170 ) );
  OR4_X1 u1_u4_u0_U72 (.ZN( u1_out4_31 ) , .A4( u1_u4_u0_n155 ) , .A2( u1_u4_u0_n156 ) , .A1( u1_u4_u0_n157 ) , .A3( u1_u4_u0_n173 ) );
  AOI21_X1 u1_u4_u0_U73 (.A( u1_u4_u0_n138 ) , .B2( u1_u4_u0_n139 ) , .B1( u1_u4_u0_n140 ) , .ZN( u1_u4_u0_n157 ) );
  AOI21_X1 u1_u4_u0_U74 (.B2( u1_u4_u0_n141 ) , .B1( u1_u4_u0_n142 ) , .ZN( u1_u4_u0_n156 ) , .A( u1_u4_u0_n161 ) );
  INV_X1 u1_u4_u0_U75 (.ZN( u1_u4_u0_n174 ) , .A( u1_u4_u0_n89 ) );
  AOI211_X1 u1_u4_u0_U76 (.B( u1_u4_u0_n104 ) , .A( u1_u4_u0_n105 ) , .ZN( u1_u4_u0_n106 ) , .C2( u1_u4_u0_n113 ) , .C1( u1_u4_u0_n160 ) );
  OR4_X1 u1_u4_u0_U77 (.ZN( u1_out4_17 ) , .A4( u1_u4_u0_n122 ) , .A2( u1_u4_u0_n123 ) , .A1( u1_u4_u0_n124 ) , .A3( u1_u4_u0_n170 ) );
  OAI221_X1 u1_u4_u0_U78 (.C1( u1_u4_u0_n121 ) , .ZN( u1_u4_u0_n122 ) , .B2( u1_u4_u0_n127 ) , .A( u1_u4_u0_n143 ) , .B1( u1_u4_u0_n144 ) , .C2( u1_u4_u0_n147 ) );
  NOR2_X1 u1_u4_u0_U79 (.A1( u1_u4_u0_n120 ) , .ZN( u1_u4_u0_n143 ) , .A2( u1_u4_u0_n167 ) );
  AND2_X1 u1_u4_u0_U8 (.A1( u1_u4_u0_n114 ) , .A2( u1_u4_u0_n121 ) , .ZN( u1_u4_u0_n146 ) );
  AOI21_X1 u1_u4_u0_U80 (.B1( u1_u4_u0_n132 ) , .ZN( u1_u4_u0_n133 ) , .A( u1_u4_u0_n144 ) , .B2( u1_u4_u0_n166 ) );
  OAI22_X1 u1_u4_u0_U81 (.ZN( u1_u4_u0_n105 ) , .A2( u1_u4_u0_n132 ) , .B1( u1_u4_u0_n146 ) , .A1( u1_u4_u0_n147 ) , .B2( u1_u4_u0_n161 ) );
  NAND2_X1 u1_u4_u0_U82 (.ZN( u1_u4_u0_n110 ) , .A2( u1_u4_u0_n132 ) , .A1( u1_u4_u0_n145 ) );
  INV_X1 u1_u4_u0_U83 (.A( u1_u4_u0_n119 ) , .ZN( u1_u4_u0_n167 ) );
  NAND2_X1 u1_u4_u0_U84 (.A2( u1_u4_u0_n103 ) , .ZN( u1_u4_u0_n140 ) , .A1( u1_u4_u0_n94 ) );
  NAND2_X1 u1_u4_u0_U85 (.A1( u1_u4_u0_n101 ) , .ZN( u1_u4_u0_n130 ) , .A2( u1_u4_u0_n94 ) );
  NAND2_X1 u1_u4_u0_U86 (.ZN( u1_u4_u0_n108 ) , .A1( u1_u4_u0_n92 ) , .A2( u1_u4_u0_n94 ) );
  NAND2_X1 u1_u4_u0_U87 (.ZN( u1_u4_u0_n142 ) , .A1( u1_u4_u0_n94 ) , .A2( u1_u4_u0_n95 ) );
  NAND3_X1 u1_u4_u0_U88 (.ZN( u1_out4_23 ) , .A3( u1_u4_u0_n137 ) , .A1( u1_u4_u0_n168 ) , .A2( u1_u4_u0_n171 ) );
  NAND3_X1 u1_u4_u0_U89 (.A3( u1_u4_u0_n127 ) , .A2( u1_u4_u0_n128 ) , .ZN( u1_u4_u0_n135 ) , .A1( u1_u4_u0_n150 ) );
  AND2_X1 u1_u4_u0_U9 (.A1( u1_u4_u0_n131 ) , .ZN( u1_u4_u0_n141 ) , .A2( u1_u4_u0_n150 ) );
  NAND3_X1 u1_u4_u0_U90 (.ZN( u1_u4_u0_n117 ) , .A3( u1_u4_u0_n132 ) , .A2( u1_u4_u0_n139 ) , .A1( u1_u4_u0_n148 ) );
  NAND3_X1 u1_u4_u0_U91 (.ZN( u1_u4_u0_n109 ) , .A2( u1_u4_u0_n114 ) , .A3( u1_u4_u0_n140 ) , .A1( u1_u4_u0_n149 ) );
  NAND3_X1 u1_u4_u0_U92 (.ZN( u1_out4_9 ) , .A3( u1_u4_u0_n106 ) , .A2( u1_u4_u0_n171 ) , .A1( u1_u4_u0_n174 ) );
  NAND3_X1 u1_u4_u0_U93 (.A2( u1_u4_u0_n128 ) , .A1( u1_u4_u0_n132 ) , .A3( u1_u4_u0_n146 ) , .ZN( u1_u4_u0_n97 ) );
  OAI22_X1 u1_u4_u2_U10 (.ZN( u1_u4_u2_n109 ) , .A2( u1_u4_u2_n113 ) , .B2( u1_u4_u2_n133 ) , .B1( u1_u4_u2_n167 ) , .A1( u1_u4_u2_n168 ) );
  NAND3_X1 u1_u4_u2_U100 (.A2( u1_u4_u2_n100 ) , .A1( u1_u4_u2_n104 ) , .A3( u1_u4_u2_n138 ) , .ZN( u1_u4_u2_n98 ) );
  OAI22_X1 u1_u4_u2_U11 (.B1( u1_u4_u2_n151 ) , .A2( u1_u4_u2_n152 ) , .A1( u1_u4_u2_n153 ) , .ZN( u1_u4_u2_n160 ) , .B2( u1_u4_u2_n168 ) );
  NOR3_X1 u1_u4_u2_U12 (.A1( u1_u4_u2_n150 ) , .ZN( u1_u4_u2_n151 ) , .A3( u1_u4_u2_n175 ) , .A2( u1_u4_u2_n188 ) );
  AOI21_X1 u1_u4_u2_U13 (.ZN( u1_u4_u2_n144 ) , .B2( u1_u4_u2_n155 ) , .A( u1_u4_u2_n172 ) , .B1( u1_u4_u2_n185 ) );
  AOI21_X1 u1_u4_u2_U14 (.B2( u1_u4_u2_n143 ) , .ZN( u1_u4_u2_n145 ) , .B1( u1_u4_u2_n152 ) , .A( u1_u4_u2_n171 ) );
  AOI21_X1 u1_u4_u2_U15 (.B2( u1_u4_u2_n120 ) , .B1( u1_u4_u2_n121 ) , .ZN( u1_u4_u2_n126 ) , .A( u1_u4_u2_n167 ) );
  INV_X1 u1_u4_u2_U16 (.A( u1_u4_u2_n156 ) , .ZN( u1_u4_u2_n171 ) );
  INV_X1 u1_u4_u2_U17 (.A( u1_u4_u2_n120 ) , .ZN( u1_u4_u2_n188 ) );
  NAND2_X1 u1_u4_u2_U18 (.A2( u1_u4_u2_n122 ) , .ZN( u1_u4_u2_n150 ) , .A1( u1_u4_u2_n152 ) );
  INV_X1 u1_u4_u2_U19 (.A( u1_u4_u2_n153 ) , .ZN( u1_u4_u2_n170 ) );
  INV_X1 u1_u4_u2_U20 (.A( u1_u4_u2_n137 ) , .ZN( u1_u4_u2_n173 ) );
  NAND2_X1 u1_u4_u2_U21 (.A1( u1_u4_u2_n132 ) , .A2( u1_u4_u2_n139 ) , .ZN( u1_u4_u2_n157 ) );
  INV_X1 u1_u4_u2_U22 (.A( u1_u4_u2_n113 ) , .ZN( u1_u4_u2_n178 ) );
  INV_X1 u1_u4_u2_U23 (.A( u1_u4_u2_n139 ) , .ZN( u1_u4_u2_n175 ) );
  INV_X1 u1_u4_u2_U24 (.A( u1_u4_u2_n155 ) , .ZN( u1_u4_u2_n181 ) );
  INV_X1 u1_u4_u2_U25 (.A( u1_u4_u2_n119 ) , .ZN( u1_u4_u2_n177 ) );
  INV_X1 u1_u4_u2_U26 (.A( u1_u4_u2_n116 ) , .ZN( u1_u4_u2_n180 ) );
  INV_X1 u1_u4_u2_U27 (.A( u1_u4_u2_n131 ) , .ZN( u1_u4_u2_n179 ) );
  INV_X1 u1_u4_u2_U28 (.A( u1_u4_u2_n154 ) , .ZN( u1_u4_u2_n176 ) );
  NAND2_X1 u1_u4_u2_U29 (.A2( u1_u4_u2_n116 ) , .A1( u1_u4_u2_n117 ) , .ZN( u1_u4_u2_n118 ) );
  NOR2_X1 u1_u4_u2_U3 (.ZN( u1_u4_u2_n121 ) , .A2( u1_u4_u2_n177 ) , .A1( u1_u4_u2_n180 ) );
  INV_X1 u1_u4_u2_U30 (.A( u1_u4_u2_n132 ) , .ZN( u1_u4_u2_n182 ) );
  INV_X1 u1_u4_u2_U31 (.A( u1_u4_u2_n158 ) , .ZN( u1_u4_u2_n183 ) );
  OAI21_X1 u1_u4_u2_U32 (.A( u1_u4_u2_n156 ) , .B1( u1_u4_u2_n157 ) , .ZN( u1_u4_u2_n158 ) , .B2( u1_u4_u2_n179 ) );
  NOR2_X1 u1_u4_u2_U33 (.ZN( u1_u4_u2_n156 ) , .A1( u1_u4_u2_n166 ) , .A2( u1_u4_u2_n169 ) );
  NOR2_X1 u1_u4_u2_U34 (.A2( u1_u4_u2_n114 ) , .ZN( u1_u4_u2_n137 ) , .A1( u1_u4_u2_n140 ) );
  NOR2_X1 u1_u4_u2_U35 (.A2( u1_u4_u2_n138 ) , .ZN( u1_u4_u2_n153 ) , .A1( u1_u4_u2_n156 ) );
  AOI211_X1 u1_u4_u2_U36 (.ZN( u1_u4_u2_n130 ) , .C1( u1_u4_u2_n138 ) , .C2( u1_u4_u2_n179 ) , .B( u1_u4_u2_n96 ) , .A( u1_u4_u2_n97 ) );
  OAI22_X1 u1_u4_u2_U37 (.B1( u1_u4_u2_n133 ) , .A2( u1_u4_u2_n137 ) , .A1( u1_u4_u2_n152 ) , .B2( u1_u4_u2_n168 ) , .ZN( u1_u4_u2_n97 ) );
  OAI221_X1 u1_u4_u2_U38 (.B1( u1_u4_u2_n113 ) , .C1( u1_u4_u2_n132 ) , .A( u1_u4_u2_n149 ) , .B2( u1_u4_u2_n171 ) , .C2( u1_u4_u2_n172 ) , .ZN( u1_u4_u2_n96 ) );
  OAI221_X1 u1_u4_u2_U39 (.A( u1_u4_u2_n115 ) , .C2( u1_u4_u2_n123 ) , .B2( u1_u4_u2_n143 ) , .B1( u1_u4_u2_n153 ) , .ZN( u1_u4_u2_n163 ) , .C1( u1_u4_u2_n168 ) );
  INV_X1 u1_u4_u2_U4 (.A( u1_u4_u2_n134 ) , .ZN( u1_u4_u2_n185 ) );
  OAI21_X1 u1_u4_u2_U40 (.A( u1_u4_u2_n114 ) , .ZN( u1_u4_u2_n115 ) , .B1( u1_u4_u2_n176 ) , .B2( u1_u4_u2_n178 ) );
  OAI221_X1 u1_u4_u2_U41 (.A( u1_u4_u2_n135 ) , .B2( u1_u4_u2_n136 ) , .B1( u1_u4_u2_n137 ) , .ZN( u1_u4_u2_n162 ) , .C2( u1_u4_u2_n167 ) , .C1( u1_u4_u2_n185 ) );
  AND3_X1 u1_u4_u2_U42 (.A3( u1_u4_u2_n131 ) , .A2( u1_u4_u2_n132 ) , .A1( u1_u4_u2_n133 ) , .ZN( u1_u4_u2_n136 ) );
  AOI22_X1 u1_u4_u2_U43 (.ZN( u1_u4_u2_n135 ) , .B1( u1_u4_u2_n140 ) , .A1( u1_u4_u2_n156 ) , .B2( u1_u4_u2_n180 ) , .A2( u1_u4_u2_n188 ) );
  AOI21_X1 u1_u4_u2_U44 (.ZN( u1_u4_u2_n149 ) , .B1( u1_u4_u2_n173 ) , .B2( u1_u4_u2_n188 ) , .A( u1_u4_u2_n95 ) );
  AND3_X1 u1_u4_u2_U45 (.A2( u1_u4_u2_n100 ) , .A1( u1_u4_u2_n104 ) , .A3( u1_u4_u2_n156 ) , .ZN( u1_u4_u2_n95 ) );
  OAI21_X1 u1_u4_u2_U46 (.A( u1_u4_u2_n101 ) , .B2( u1_u4_u2_n121 ) , .B1( u1_u4_u2_n153 ) , .ZN( u1_u4_u2_n164 ) );
  NAND2_X1 u1_u4_u2_U47 (.A2( u1_u4_u2_n100 ) , .A1( u1_u4_u2_n107 ) , .ZN( u1_u4_u2_n155 ) );
  NAND2_X1 u1_u4_u2_U48 (.A2( u1_u4_u2_n105 ) , .A1( u1_u4_u2_n108 ) , .ZN( u1_u4_u2_n143 ) );
  NAND2_X1 u1_u4_u2_U49 (.A1( u1_u4_u2_n104 ) , .A2( u1_u4_u2_n106 ) , .ZN( u1_u4_u2_n152 ) );
  INV_X1 u1_u4_u2_U5 (.A( u1_u4_u2_n150 ) , .ZN( u1_u4_u2_n184 ) );
  NAND2_X1 u1_u4_u2_U50 (.A1( u1_u4_u2_n100 ) , .A2( u1_u4_u2_n105 ) , .ZN( u1_u4_u2_n132 ) );
  INV_X1 u1_u4_u2_U51 (.A( u1_u4_u2_n140 ) , .ZN( u1_u4_u2_n168 ) );
  INV_X1 u1_u4_u2_U52 (.A( u1_u4_u2_n138 ) , .ZN( u1_u4_u2_n167 ) );
  OAI21_X1 u1_u4_u2_U53 (.A( u1_u4_u2_n141 ) , .B2( u1_u4_u2_n142 ) , .ZN( u1_u4_u2_n146 ) , .B1( u1_u4_u2_n153 ) );
  OAI21_X1 u1_u4_u2_U54 (.A( u1_u4_u2_n140 ) , .ZN( u1_u4_u2_n141 ) , .B1( u1_u4_u2_n176 ) , .B2( u1_u4_u2_n177 ) );
  NOR3_X1 u1_u4_u2_U55 (.ZN( u1_u4_u2_n142 ) , .A3( u1_u4_u2_n175 ) , .A2( u1_u4_u2_n178 ) , .A1( u1_u4_u2_n181 ) );
  INV_X1 u1_u4_u2_U56 (.ZN( u1_u4_u2_n187 ) , .A( u1_u4_u2_n99 ) );
  OAI21_X1 u1_u4_u2_U57 (.B1( u1_u4_u2_n137 ) , .B2( u1_u4_u2_n143 ) , .A( u1_u4_u2_n98 ) , .ZN( u1_u4_u2_n99 ) );
  NAND2_X1 u1_u4_u2_U58 (.A1( u1_u4_u2_n102 ) , .A2( u1_u4_u2_n106 ) , .ZN( u1_u4_u2_n113 ) );
  NAND2_X1 u1_u4_u2_U59 (.A1( u1_u4_u2_n106 ) , .A2( u1_u4_u2_n107 ) , .ZN( u1_u4_u2_n131 ) );
  NOR4_X1 u1_u4_u2_U6 (.A4( u1_u4_u2_n124 ) , .A3( u1_u4_u2_n125 ) , .A2( u1_u4_u2_n126 ) , .A1( u1_u4_u2_n127 ) , .ZN( u1_u4_u2_n128 ) );
  NAND2_X1 u1_u4_u2_U60 (.A1( u1_u4_u2_n103 ) , .A2( u1_u4_u2_n107 ) , .ZN( u1_u4_u2_n139 ) );
  NAND2_X1 u1_u4_u2_U61 (.A1( u1_u4_u2_n103 ) , .A2( u1_u4_u2_n105 ) , .ZN( u1_u4_u2_n133 ) );
  NAND2_X1 u1_u4_u2_U62 (.A1( u1_u4_u2_n102 ) , .A2( u1_u4_u2_n103 ) , .ZN( u1_u4_u2_n154 ) );
  NAND2_X1 u1_u4_u2_U63 (.A2( u1_u4_u2_n103 ) , .A1( u1_u4_u2_n104 ) , .ZN( u1_u4_u2_n119 ) );
  NAND2_X1 u1_u4_u2_U64 (.A2( u1_u4_u2_n107 ) , .A1( u1_u4_u2_n108 ) , .ZN( u1_u4_u2_n123 ) );
  NAND2_X1 u1_u4_u2_U65 (.A1( u1_u4_u2_n104 ) , .A2( u1_u4_u2_n108 ) , .ZN( u1_u4_u2_n122 ) );
  INV_X1 u1_u4_u2_U66 (.A( u1_u4_u2_n114 ) , .ZN( u1_u4_u2_n172 ) );
  NAND2_X1 u1_u4_u2_U67 (.A2( u1_u4_u2_n100 ) , .A1( u1_u4_u2_n102 ) , .ZN( u1_u4_u2_n116 ) );
  NAND2_X1 u1_u4_u2_U68 (.A1( u1_u4_u2_n102 ) , .A2( u1_u4_u2_n108 ) , .ZN( u1_u4_u2_n120 ) );
  NAND2_X1 u1_u4_u2_U69 (.A2( u1_u4_u2_n105 ) , .A1( u1_u4_u2_n106 ) , .ZN( u1_u4_u2_n117 ) );
  AOI21_X1 u1_u4_u2_U7 (.B2( u1_u4_u2_n119 ) , .ZN( u1_u4_u2_n127 ) , .A( u1_u4_u2_n137 ) , .B1( u1_u4_u2_n155 ) );
  NOR2_X1 u1_u4_u2_U70 (.A2( u1_u4_X_16 ) , .ZN( u1_u4_u2_n140 ) , .A1( u1_u4_u2_n166 ) );
  NOR2_X1 u1_u4_u2_U71 (.A2( u1_u4_X_13 ) , .A1( u1_u4_X_14 ) , .ZN( u1_u4_u2_n100 ) );
  NOR2_X1 u1_u4_u2_U72 (.A2( u1_u4_X_16 ) , .A1( u1_u4_X_17 ) , .ZN( u1_u4_u2_n138 ) );
  NOR2_X1 u1_u4_u2_U73 (.A2( u1_u4_X_15 ) , .A1( u1_u4_X_18 ) , .ZN( u1_u4_u2_n104 ) );
  NOR2_X1 u1_u4_u2_U74 (.A2( u1_u4_X_14 ) , .ZN( u1_u4_u2_n103 ) , .A1( u1_u4_u2_n174 ) );
  NOR2_X1 u1_u4_u2_U75 (.A2( u1_u4_X_15 ) , .ZN( u1_u4_u2_n102 ) , .A1( u1_u4_u2_n165 ) );
  NOR2_X1 u1_u4_u2_U76 (.A2( u1_u4_X_17 ) , .ZN( u1_u4_u2_n114 ) , .A1( u1_u4_u2_n169 ) );
  AND2_X1 u1_u4_u2_U77 (.A1( u1_u4_X_15 ) , .ZN( u1_u4_u2_n105 ) , .A2( u1_u4_u2_n165 ) );
  AND2_X1 u1_u4_u2_U78 (.A2( u1_u4_X_15 ) , .A1( u1_u4_X_18 ) , .ZN( u1_u4_u2_n107 ) );
  AND2_X1 u1_u4_u2_U79 (.A1( u1_u4_X_14 ) , .ZN( u1_u4_u2_n106 ) , .A2( u1_u4_u2_n174 ) );
  AOI21_X1 u1_u4_u2_U8 (.ZN( u1_u4_u2_n124 ) , .B1( u1_u4_u2_n131 ) , .B2( u1_u4_u2_n143 ) , .A( u1_u4_u2_n172 ) );
  AND2_X1 u1_u4_u2_U80 (.A1( u1_u4_X_13 ) , .A2( u1_u4_X_14 ) , .ZN( u1_u4_u2_n108 ) );
  INV_X1 u1_u4_u2_U81 (.A( u1_u4_X_16 ) , .ZN( u1_u4_u2_n169 ) );
  INV_X1 u1_u4_u2_U82 (.A( u1_u4_X_17 ) , .ZN( u1_u4_u2_n166 ) );
  INV_X1 u1_u4_u2_U83 (.A( u1_u4_X_13 ) , .ZN( u1_u4_u2_n174 ) );
  INV_X1 u1_u4_u2_U84 (.A( u1_u4_X_18 ) , .ZN( u1_u4_u2_n165 ) );
  NAND4_X1 u1_u4_u2_U85 (.ZN( u1_out4_30 ) , .A4( u1_u4_u2_n147 ) , .A3( u1_u4_u2_n148 ) , .A2( u1_u4_u2_n149 ) , .A1( u1_u4_u2_n187 ) );
  NOR3_X1 u1_u4_u2_U86 (.A3( u1_u4_u2_n144 ) , .A2( u1_u4_u2_n145 ) , .A1( u1_u4_u2_n146 ) , .ZN( u1_u4_u2_n147 ) );
  AOI21_X1 u1_u4_u2_U87 (.B2( u1_u4_u2_n138 ) , .ZN( u1_u4_u2_n148 ) , .A( u1_u4_u2_n162 ) , .B1( u1_u4_u2_n182 ) );
  NAND4_X1 u1_u4_u2_U88 (.ZN( u1_out4_24 ) , .A4( u1_u4_u2_n111 ) , .A3( u1_u4_u2_n112 ) , .A1( u1_u4_u2_n130 ) , .A2( u1_u4_u2_n187 ) );
  AOI221_X1 u1_u4_u2_U89 (.A( u1_u4_u2_n109 ) , .B1( u1_u4_u2_n110 ) , .ZN( u1_u4_u2_n111 ) , .C1( u1_u4_u2_n134 ) , .C2( u1_u4_u2_n170 ) , .B2( u1_u4_u2_n173 ) );
  AOI21_X1 u1_u4_u2_U9 (.B2( u1_u4_u2_n123 ) , .ZN( u1_u4_u2_n125 ) , .A( u1_u4_u2_n171 ) , .B1( u1_u4_u2_n184 ) );
  AOI21_X1 u1_u4_u2_U90 (.ZN( u1_u4_u2_n112 ) , .B2( u1_u4_u2_n156 ) , .A( u1_u4_u2_n164 ) , .B1( u1_u4_u2_n181 ) );
  NAND4_X1 u1_u4_u2_U91 (.ZN( u1_out4_16 ) , .A4( u1_u4_u2_n128 ) , .A3( u1_u4_u2_n129 ) , .A1( u1_u4_u2_n130 ) , .A2( u1_u4_u2_n186 ) );
  AOI22_X1 u1_u4_u2_U92 (.A2( u1_u4_u2_n118 ) , .ZN( u1_u4_u2_n129 ) , .A1( u1_u4_u2_n140 ) , .B1( u1_u4_u2_n157 ) , .B2( u1_u4_u2_n170 ) );
  INV_X1 u1_u4_u2_U93 (.A( u1_u4_u2_n163 ) , .ZN( u1_u4_u2_n186 ) );
  OR4_X1 u1_u4_u2_U94 (.ZN( u1_out4_6 ) , .A4( u1_u4_u2_n161 ) , .A3( u1_u4_u2_n162 ) , .A2( u1_u4_u2_n163 ) , .A1( u1_u4_u2_n164 ) );
  OR3_X1 u1_u4_u2_U95 (.A2( u1_u4_u2_n159 ) , .A1( u1_u4_u2_n160 ) , .ZN( u1_u4_u2_n161 ) , .A3( u1_u4_u2_n183 ) );
  AOI21_X1 u1_u4_u2_U96 (.B2( u1_u4_u2_n154 ) , .B1( u1_u4_u2_n155 ) , .ZN( u1_u4_u2_n159 ) , .A( u1_u4_u2_n167 ) );
  NAND3_X1 u1_u4_u2_U97 (.A2( u1_u4_u2_n117 ) , .A1( u1_u4_u2_n122 ) , .A3( u1_u4_u2_n123 ) , .ZN( u1_u4_u2_n134 ) );
  NAND3_X1 u1_u4_u2_U98 (.ZN( u1_u4_u2_n110 ) , .A2( u1_u4_u2_n131 ) , .A3( u1_u4_u2_n139 ) , .A1( u1_u4_u2_n154 ) );
  NAND3_X1 u1_u4_u2_U99 (.A2( u1_u4_u2_n100 ) , .ZN( u1_u4_u2_n101 ) , .A1( u1_u4_u2_n104 ) , .A3( u1_u4_u2_n114 ) );
  XOR2_X1 u1_u6_U16 (.B( u1_K7_3 ) , .A( u1_R5_2 ) , .Z( u1_u6_X_3 ) );
  XOR2_X1 u1_u6_U20 (.B( u1_K7_36 ) , .A( u1_R5_25 ) , .Z( u1_u6_X_36 ) );
  XOR2_X1 u1_u6_U21 (.B( u1_K7_35 ) , .A( u1_R5_24 ) , .Z( u1_u6_X_35 ) );
  XOR2_X1 u1_u6_U22 (.B( u1_K7_34 ) , .A( u1_R5_23 ) , .Z( u1_u6_X_34 ) );
  XOR2_X1 u1_u6_U23 (.B( u1_K7_33 ) , .A( u1_R5_22 ) , .Z( u1_u6_X_33 ) );
  XOR2_X1 u1_u6_U24 (.B( u1_K7_32 ) , .A( u1_R5_21 ) , .Z( u1_u6_X_32 ) );
  XOR2_X1 u1_u6_U25 (.B( u1_K7_31 ) , .A( u1_R5_20 ) , .Z( u1_u6_X_31 ) );
  XOR2_X1 u1_u6_U27 (.B( u1_K7_2 ) , .A( u1_R5_1 ) , .Z( u1_u6_X_2 ) );
  XOR2_X1 u1_u6_U38 (.B( u1_K7_1 ) , .A( u1_R5_32 ) , .Z( u1_u6_X_1 ) );
  XOR2_X1 u1_u6_U4 (.B( u1_K7_6 ) , .A( u1_R5_5 ) , .Z( u1_u6_X_6 ) );
  XOR2_X1 u1_u6_U5 (.B( u1_K7_5 ) , .A( u1_R5_4 ) , .Z( u1_u6_X_5 ) );
  XOR2_X1 u1_u6_U6 (.B( u1_K7_4 ) , .A( u1_R5_3 ) , .Z( u1_u6_X_4 ) );
  AND3_X1 u1_u6_u0_U10 (.A2( u1_u6_u0_n112 ) , .ZN( u1_u6_u0_n127 ) , .A3( u1_u6_u0_n130 ) , .A1( u1_u6_u0_n148 ) );
  NAND2_X1 u1_u6_u0_U11 (.ZN( u1_u6_u0_n113 ) , .A1( u1_u6_u0_n139 ) , .A2( u1_u6_u0_n149 ) );
  AND2_X1 u1_u6_u0_U12 (.ZN( u1_u6_u0_n107 ) , .A1( u1_u6_u0_n130 ) , .A2( u1_u6_u0_n140 ) );
  AND2_X1 u1_u6_u0_U13 (.A2( u1_u6_u0_n129 ) , .A1( u1_u6_u0_n130 ) , .ZN( u1_u6_u0_n151 ) );
  AND2_X1 u1_u6_u0_U14 (.A1( u1_u6_u0_n108 ) , .A2( u1_u6_u0_n125 ) , .ZN( u1_u6_u0_n145 ) );
  INV_X1 u1_u6_u0_U15 (.A( u1_u6_u0_n143 ) , .ZN( u1_u6_u0_n173 ) );
  NOR2_X1 u1_u6_u0_U16 (.A2( u1_u6_u0_n136 ) , .ZN( u1_u6_u0_n147 ) , .A1( u1_u6_u0_n160 ) );
  NOR2_X1 u1_u6_u0_U17 (.A1( u1_u6_u0_n163 ) , .A2( u1_u6_u0_n164 ) , .ZN( u1_u6_u0_n95 ) );
  AOI21_X1 u1_u6_u0_U18 (.B1( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n132 ) , .A( u1_u6_u0_n165 ) , .B2( u1_u6_u0_n93 ) );
  INV_X1 u1_u6_u0_U19 (.A( u1_u6_u0_n142 ) , .ZN( u1_u6_u0_n165 ) );
  OAI221_X1 u1_u6_u0_U20 (.C1( u1_u6_u0_n112 ) , .ZN( u1_u6_u0_n120 ) , .B1( u1_u6_u0_n138 ) , .B2( u1_u6_u0_n141 ) , .C2( u1_u6_u0_n147 ) , .A( u1_u6_u0_n172 ) );
  AOI211_X1 u1_u6_u0_U21 (.B( u1_u6_u0_n115 ) , .A( u1_u6_u0_n116 ) , .C2( u1_u6_u0_n117 ) , .C1( u1_u6_u0_n118 ) , .ZN( u1_u6_u0_n119 ) );
  OAI22_X1 u1_u6_u0_U22 (.B1( u1_u6_u0_n125 ) , .ZN( u1_u6_u0_n126 ) , .A1( u1_u6_u0_n138 ) , .A2( u1_u6_u0_n146 ) , .B2( u1_u6_u0_n147 ) );
  OAI22_X1 u1_u6_u0_U23 (.B1( u1_u6_u0_n131 ) , .A1( u1_u6_u0_n144 ) , .B2( u1_u6_u0_n147 ) , .A2( u1_u6_u0_n90 ) , .ZN( u1_u6_u0_n91 ) );
  AND3_X1 u1_u6_u0_U24 (.A3( u1_u6_u0_n121 ) , .A2( u1_u6_u0_n125 ) , .A1( u1_u6_u0_n148 ) , .ZN( u1_u6_u0_n90 ) );
  NAND2_X1 u1_u6_u0_U25 (.A1( u1_u6_u0_n100 ) , .A2( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n125 ) );
  INV_X1 u1_u6_u0_U26 (.A( u1_u6_u0_n136 ) , .ZN( u1_u6_u0_n161 ) );
  AOI22_X1 u1_u6_u0_U27 (.B2( u1_u6_u0_n109 ) , .A2( u1_u6_u0_n110 ) , .ZN( u1_u6_u0_n111 ) , .B1( u1_u6_u0_n118 ) , .A1( u1_u6_u0_n160 ) );
  NAND2_X1 u1_u6_u0_U28 (.A1( u1_u6_u0_n100 ) , .ZN( u1_u6_u0_n129 ) , .A2( u1_u6_u0_n95 ) );
  INV_X1 u1_u6_u0_U29 (.A( u1_u6_u0_n118 ) , .ZN( u1_u6_u0_n158 ) );
  INV_X1 u1_u6_u0_U3 (.A( u1_u6_u0_n113 ) , .ZN( u1_u6_u0_n166 ) );
  AOI21_X1 u1_u6_u0_U30 (.ZN( u1_u6_u0_n104 ) , .B1( u1_u6_u0_n107 ) , .B2( u1_u6_u0_n141 ) , .A( u1_u6_u0_n144 ) );
  AOI21_X1 u1_u6_u0_U31 (.B1( u1_u6_u0_n127 ) , .B2( u1_u6_u0_n129 ) , .A( u1_u6_u0_n138 ) , .ZN( u1_u6_u0_n96 ) );
  AOI21_X1 u1_u6_u0_U32 (.ZN( u1_u6_u0_n116 ) , .B2( u1_u6_u0_n142 ) , .A( u1_u6_u0_n144 ) , .B1( u1_u6_u0_n166 ) );
  NAND2_X1 u1_u6_u0_U33 (.A2( u1_u6_u0_n100 ) , .A1( u1_u6_u0_n101 ) , .ZN( u1_u6_u0_n139 ) );
  NAND2_X1 u1_u6_u0_U34 (.A2( u1_u6_u0_n100 ) , .ZN( u1_u6_u0_n131 ) , .A1( u1_u6_u0_n92 ) );
  NAND2_X1 u1_u6_u0_U35 (.A1( u1_u6_u0_n101 ) , .A2( u1_u6_u0_n102 ) , .ZN( u1_u6_u0_n150 ) );
  INV_X1 u1_u6_u0_U36 (.A( u1_u6_u0_n138 ) , .ZN( u1_u6_u0_n160 ) );
  NAND2_X1 u1_u6_u0_U37 (.A1( u1_u6_u0_n102 ) , .ZN( u1_u6_u0_n128 ) , .A2( u1_u6_u0_n95 ) );
  NAND2_X1 u1_u6_u0_U38 (.ZN( u1_u6_u0_n148 ) , .A1( u1_u6_u0_n93 ) , .A2( u1_u6_u0_n95 ) );
  NAND2_X1 u1_u6_u0_U39 (.A2( u1_u6_u0_n102 ) , .A1( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n149 ) );
  AOI21_X1 u1_u6_u0_U4 (.B1( u1_u6_u0_n114 ) , .ZN( u1_u6_u0_n115 ) , .B2( u1_u6_u0_n129 ) , .A( u1_u6_u0_n161 ) );
  NAND2_X1 u1_u6_u0_U40 (.A2( u1_u6_u0_n102 ) , .ZN( u1_u6_u0_n114 ) , .A1( u1_u6_u0_n92 ) );
  NAND2_X1 u1_u6_u0_U41 (.A2( u1_u6_u0_n101 ) , .ZN( u1_u6_u0_n121 ) , .A1( u1_u6_u0_n93 ) );
  NAND2_X1 u1_u6_u0_U42 (.ZN( u1_u6_u0_n112 ) , .A2( u1_u6_u0_n92 ) , .A1( u1_u6_u0_n93 ) );
  INV_X1 u1_u6_u0_U43 (.ZN( u1_u6_u0_n172 ) , .A( u1_u6_u0_n88 ) );
  OAI222_X1 u1_u6_u0_U44 (.C1( u1_u6_u0_n108 ) , .A1( u1_u6_u0_n125 ) , .B2( u1_u6_u0_n128 ) , .B1( u1_u6_u0_n144 ) , .A2( u1_u6_u0_n158 ) , .C2( u1_u6_u0_n161 ) , .ZN( u1_u6_u0_n88 ) );
  OR3_X1 u1_u6_u0_U45 (.A3( u1_u6_u0_n152 ) , .A2( u1_u6_u0_n153 ) , .A1( u1_u6_u0_n154 ) , .ZN( u1_u6_u0_n155 ) );
  AOI21_X1 u1_u6_u0_U46 (.A( u1_u6_u0_n144 ) , .B2( u1_u6_u0_n145 ) , .B1( u1_u6_u0_n146 ) , .ZN( u1_u6_u0_n154 ) );
  AOI21_X1 u1_u6_u0_U47 (.B2( u1_u6_u0_n150 ) , .B1( u1_u6_u0_n151 ) , .ZN( u1_u6_u0_n152 ) , .A( u1_u6_u0_n158 ) );
  AOI21_X1 u1_u6_u0_U48 (.A( u1_u6_u0_n147 ) , .B2( u1_u6_u0_n148 ) , .B1( u1_u6_u0_n149 ) , .ZN( u1_u6_u0_n153 ) );
  INV_X1 u1_u6_u0_U49 (.ZN( u1_u6_u0_n171 ) , .A( u1_u6_u0_n99 ) );
  AOI21_X1 u1_u6_u0_U5 (.B2( u1_u6_u0_n131 ) , .ZN( u1_u6_u0_n134 ) , .B1( u1_u6_u0_n151 ) , .A( u1_u6_u0_n158 ) );
  OAI211_X1 u1_u6_u0_U50 (.C2( u1_u6_u0_n140 ) , .C1( u1_u6_u0_n161 ) , .A( u1_u6_u0_n169 ) , .B( u1_u6_u0_n98 ) , .ZN( u1_u6_u0_n99 ) );
  INV_X1 u1_u6_u0_U51 (.ZN( u1_u6_u0_n169 ) , .A( u1_u6_u0_n91 ) );
  AOI211_X1 u1_u6_u0_U52 (.C1( u1_u6_u0_n118 ) , .A( u1_u6_u0_n123 ) , .B( u1_u6_u0_n96 ) , .C2( u1_u6_u0_n97 ) , .ZN( u1_u6_u0_n98 ) );
  NOR2_X1 u1_u6_u0_U53 (.A2( u1_u6_X_4 ) , .A1( u1_u6_X_5 ) , .ZN( u1_u6_u0_n118 ) );
  NOR2_X1 u1_u6_u0_U54 (.A2( u1_u6_X_2 ) , .ZN( u1_u6_u0_n103 ) , .A1( u1_u6_u0_n164 ) );
  NOR2_X1 u1_u6_u0_U55 (.A2( u1_u6_X_1 ) , .A1( u1_u6_X_2 ) , .ZN( u1_u6_u0_n92 ) );
  NOR2_X1 u1_u6_u0_U56 (.A2( u1_u6_X_1 ) , .ZN( u1_u6_u0_n101 ) , .A1( u1_u6_u0_n163 ) );
  NAND2_X1 u1_u6_u0_U57 (.A2( u1_u6_X_4 ) , .A1( u1_u6_X_5 ) , .ZN( u1_u6_u0_n144 ) );
  NOR2_X1 u1_u6_u0_U58 (.A2( u1_u6_X_5 ) , .ZN( u1_u6_u0_n136 ) , .A1( u1_u6_u0_n159 ) );
  NAND2_X1 u1_u6_u0_U59 (.A1( u1_u6_X_5 ) , .ZN( u1_u6_u0_n138 ) , .A2( u1_u6_u0_n159 ) );
  NOR2_X1 u1_u6_u0_U6 (.A1( u1_u6_u0_n108 ) , .ZN( u1_u6_u0_n123 ) , .A2( u1_u6_u0_n158 ) );
  AND2_X1 u1_u6_u0_U60 (.A2( u1_u6_X_3 ) , .A1( u1_u6_X_6 ) , .ZN( u1_u6_u0_n102 ) );
  INV_X1 u1_u6_u0_U61 (.A( u1_u6_X_4 ) , .ZN( u1_u6_u0_n159 ) );
  INV_X1 u1_u6_u0_U62 (.A( u1_u6_X_1 ) , .ZN( u1_u6_u0_n164 ) );
  INV_X1 u1_u6_u0_U63 (.A( u1_u6_X_2 ) , .ZN( u1_u6_u0_n163 ) );
  INV_X1 u1_u6_u0_U64 (.A( u1_u6_X_3 ) , .ZN( u1_u6_u0_n162 ) );
  INV_X1 u1_u6_u0_U65 (.A( u1_u6_u0_n126 ) , .ZN( u1_u6_u0_n168 ) );
  AOI211_X1 u1_u6_u0_U66 (.B( u1_u6_u0_n133 ) , .A( u1_u6_u0_n134 ) , .C2( u1_u6_u0_n135 ) , .C1( u1_u6_u0_n136 ) , .ZN( u1_u6_u0_n137 ) );
  OR4_X1 u1_u6_u0_U67 (.ZN( u1_out6_17 ) , .A4( u1_u6_u0_n122 ) , .A2( u1_u6_u0_n123 ) , .A1( u1_u6_u0_n124 ) , .A3( u1_u6_u0_n170 ) );
  AOI21_X1 u1_u6_u0_U68 (.B2( u1_u6_u0_n107 ) , .ZN( u1_u6_u0_n124 ) , .B1( u1_u6_u0_n128 ) , .A( u1_u6_u0_n161 ) );
  INV_X1 u1_u6_u0_U69 (.A( u1_u6_u0_n111 ) , .ZN( u1_u6_u0_n170 ) );
  OAI21_X1 u1_u6_u0_U7 (.B1( u1_u6_u0_n150 ) , .B2( u1_u6_u0_n158 ) , .A( u1_u6_u0_n172 ) , .ZN( u1_u6_u0_n89 ) );
  OR4_X1 u1_u6_u0_U70 (.ZN( u1_out6_31 ) , .A4( u1_u6_u0_n155 ) , .A2( u1_u6_u0_n156 ) , .A1( u1_u6_u0_n157 ) , .A3( u1_u6_u0_n173 ) );
  AOI21_X1 u1_u6_u0_U71 (.A( u1_u6_u0_n138 ) , .B2( u1_u6_u0_n139 ) , .B1( u1_u6_u0_n140 ) , .ZN( u1_u6_u0_n157 ) );
  AOI21_X1 u1_u6_u0_U72 (.B2( u1_u6_u0_n141 ) , .B1( u1_u6_u0_n142 ) , .ZN( u1_u6_u0_n156 ) , .A( u1_u6_u0_n161 ) );
  INV_X1 u1_u6_u0_U73 (.ZN( u1_u6_u0_n174 ) , .A( u1_u6_u0_n89 ) );
  AOI211_X1 u1_u6_u0_U74 (.B( u1_u6_u0_n104 ) , .A( u1_u6_u0_n105 ) , .ZN( u1_u6_u0_n106 ) , .C2( u1_u6_u0_n113 ) , .C1( u1_u6_u0_n160 ) );
  OAI221_X1 u1_u6_u0_U75 (.C1( u1_u6_u0_n121 ) , .ZN( u1_u6_u0_n122 ) , .B2( u1_u6_u0_n127 ) , .A( u1_u6_u0_n143 ) , .B1( u1_u6_u0_n144 ) , .C2( u1_u6_u0_n147 ) );
  NOR2_X1 u1_u6_u0_U76 (.A1( u1_u6_u0_n120 ) , .ZN( u1_u6_u0_n143 ) , .A2( u1_u6_u0_n167 ) );
  AOI21_X1 u1_u6_u0_U77 (.B1( u1_u6_u0_n132 ) , .ZN( u1_u6_u0_n133 ) , .A( u1_u6_u0_n144 ) , .B2( u1_u6_u0_n166 ) );
  OAI22_X1 u1_u6_u0_U78 (.ZN( u1_u6_u0_n105 ) , .A2( u1_u6_u0_n132 ) , .B1( u1_u6_u0_n146 ) , .A1( u1_u6_u0_n147 ) , .B2( u1_u6_u0_n161 ) );
  NAND2_X1 u1_u6_u0_U79 (.ZN( u1_u6_u0_n110 ) , .A2( u1_u6_u0_n132 ) , .A1( u1_u6_u0_n145 ) );
  AND2_X1 u1_u6_u0_U8 (.A1( u1_u6_u0_n114 ) , .A2( u1_u6_u0_n121 ) , .ZN( u1_u6_u0_n146 ) );
  INV_X1 u1_u6_u0_U80 (.A( u1_u6_u0_n119 ) , .ZN( u1_u6_u0_n167 ) );
  NAND2_X1 u1_u6_u0_U81 (.A2( u1_u6_u0_n103 ) , .ZN( u1_u6_u0_n140 ) , .A1( u1_u6_u0_n94 ) );
  NAND2_X1 u1_u6_u0_U82 (.A1( u1_u6_u0_n101 ) , .ZN( u1_u6_u0_n130 ) , .A2( u1_u6_u0_n94 ) );
  NAND2_X1 u1_u6_u0_U83 (.ZN( u1_u6_u0_n108 ) , .A1( u1_u6_u0_n92 ) , .A2( u1_u6_u0_n94 ) );
  AND2_X1 u1_u6_u0_U84 (.A1( u1_u6_X_6 ) , .A2( u1_u6_u0_n162 ) , .ZN( u1_u6_u0_n93 ) );
  NAND2_X1 u1_u6_u0_U85 (.ZN( u1_u6_u0_n142 ) , .A1( u1_u6_u0_n94 ) , .A2( u1_u6_u0_n95 ) );
  NOR2_X1 u1_u6_u0_U86 (.A2( u1_u6_X_6 ) , .ZN( u1_u6_u0_n100 ) , .A1( u1_u6_u0_n162 ) );
  NOR2_X1 u1_u6_u0_U87 (.A2( u1_u6_X_3 ) , .A1( u1_u6_X_6 ) , .ZN( u1_u6_u0_n94 ) );
  NAND3_X1 u1_u6_u0_U88 (.ZN( u1_out6_23 ) , .A3( u1_u6_u0_n137 ) , .A1( u1_u6_u0_n168 ) , .A2( u1_u6_u0_n171 ) );
  NAND3_X1 u1_u6_u0_U89 (.A3( u1_u6_u0_n127 ) , .A2( u1_u6_u0_n128 ) , .ZN( u1_u6_u0_n135 ) , .A1( u1_u6_u0_n150 ) );
  AND2_X1 u1_u6_u0_U9 (.A1( u1_u6_u0_n131 ) , .ZN( u1_u6_u0_n141 ) , .A2( u1_u6_u0_n150 ) );
  NAND3_X1 u1_u6_u0_U90 (.ZN( u1_u6_u0_n117 ) , .A3( u1_u6_u0_n132 ) , .A2( u1_u6_u0_n139 ) , .A1( u1_u6_u0_n148 ) );
  NAND3_X1 u1_u6_u0_U91 (.ZN( u1_u6_u0_n109 ) , .A2( u1_u6_u0_n114 ) , .A3( u1_u6_u0_n140 ) , .A1( u1_u6_u0_n149 ) );
  NAND3_X1 u1_u6_u0_U92 (.ZN( u1_out6_9 ) , .A3( u1_u6_u0_n106 ) , .A2( u1_u6_u0_n171 ) , .A1( u1_u6_u0_n174 ) );
  NAND3_X1 u1_u6_u0_U93 (.A2( u1_u6_u0_n128 ) , .A1( u1_u6_u0_n132 ) , .A3( u1_u6_u0_n146 ) , .ZN( u1_u6_u0_n97 ) );
  INV_X1 u1_u6_u5_U10 (.A( u1_u6_u5_n121 ) , .ZN( u1_u6_u5_n177 ) );
  AOI222_X1 u1_u6_u5_U100 (.ZN( u1_u6_u5_n113 ) , .A1( u1_u6_u5_n131 ) , .C1( u1_u6_u5_n148 ) , .B2( u1_u6_u5_n174 ) , .C2( u1_u6_u5_n178 ) , .A2( u1_u6_u5_n179 ) , .B1( u1_u6_u5_n99 ) );
  NAND4_X1 u1_u6_u5_U101 (.ZN( u1_out6_11 ) , .A4( u1_u6_u5_n143 ) , .A3( u1_u6_u5_n144 ) , .A2( u1_u6_u5_n169 ) , .A1( u1_u6_u5_n196 ) );
  AOI22_X1 u1_u6_u5_U102 (.A2( u1_u6_u5_n132 ) , .ZN( u1_u6_u5_n144 ) , .B2( u1_u6_u5_n145 ) , .B1( u1_u6_u5_n184 ) , .A1( u1_u6_u5_n194 ) );
  NOR3_X1 u1_u6_u5_U103 (.A3( u1_u6_u5_n141 ) , .A1( u1_u6_u5_n142 ) , .ZN( u1_u6_u5_n143 ) , .A2( u1_u6_u5_n191 ) );
  NAND3_X1 u1_u6_u5_U104 (.A2( u1_u6_u5_n154 ) , .A3( u1_u6_u5_n158 ) , .A1( u1_u6_u5_n161 ) , .ZN( u1_u6_u5_n99 ) );
  NOR2_X1 u1_u6_u5_U11 (.ZN( u1_u6_u5_n160 ) , .A2( u1_u6_u5_n173 ) , .A1( u1_u6_u5_n177 ) );
  INV_X1 u1_u6_u5_U12 (.A( u1_u6_u5_n150 ) , .ZN( u1_u6_u5_n174 ) );
  AOI21_X1 u1_u6_u5_U13 (.A( u1_u6_u5_n160 ) , .B2( u1_u6_u5_n161 ) , .ZN( u1_u6_u5_n162 ) , .B1( u1_u6_u5_n192 ) );
  INV_X1 u1_u6_u5_U14 (.A( u1_u6_u5_n159 ) , .ZN( u1_u6_u5_n192 ) );
  AOI21_X1 u1_u6_u5_U15 (.A( u1_u6_u5_n156 ) , .B2( u1_u6_u5_n157 ) , .B1( u1_u6_u5_n158 ) , .ZN( u1_u6_u5_n163 ) );
  AOI21_X1 u1_u6_u5_U16 (.B2( u1_u6_u5_n139 ) , .B1( u1_u6_u5_n140 ) , .ZN( u1_u6_u5_n141 ) , .A( u1_u6_u5_n150 ) );
  OAI21_X1 u1_u6_u5_U17 (.A( u1_u6_u5_n133 ) , .B2( u1_u6_u5_n134 ) , .B1( u1_u6_u5_n135 ) , .ZN( u1_u6_u5_n142 ) );
  OAI21_X1 u1_u6_u5_U18 (.ZN( u1_u6_u5_n133 ) , .B2( u1_u6_u5_n147 ) , .A( u1_u6_u5_n173 ) , .B1( u1_u6_u5_n188 ) );
  NAND2_X1 u1_u6_u5_U19 (.A2( u1_u6_u5_n119 ) , .A1( u1_u6_u5_n123 ) , .ZN( u1_u6_u5_n137 ) );
  INV_X1 u1_u6_u5_U20 (.A( u1_u6_u5_n155 ) , .ZN( u1_u6_u5_n194 ) );
  NAND2_X1 u1_u6_u5_U21 (.A1( u1_u6_u5_n121 ) , .ZN( u1_u6_u5_n132 ) , .A2( u1_u6_u5_n172 ) );
  NAND2_X1 u1_u6_u5_U22 (.A2( u1_u6_u5_n122 ) , .ZN( u1_u6_u5_n136 ) , .A1( u1_u6_u5_n154 ) );
  NAND2_X1 u1_u6_u5_U23 (.A2( u1_u6_u5_n119 ) , .A1( u1_u6_u5_n120 ) , .ZN( u1_u6_u5_n159 ) );
  INV_X1 u1_u6_u5_U24 (.A( u1_u6_u5_n156 ) , .ZN( u1_u6_u5_n175 ) );
  INV_X1 u1_u6_u5_U25 (.A( u1_u6_u5_n158 ) , .ZN( u1_u6_u5_n188 ) );
  INV_X1 u1_u6_u5_U26 (.A( u1_u6_u5_n152 ) , .ZN( u1_u6_u5_n179 ) );
  INV_X1 u1_u6_u5_U27 (.A( u1_u6_u5_n140 ) , .ZN( u1_u6_u5_n182 ) );
  INV_X1 u1_u6_u5_U28 (.A( u1_u6_u5_n151 ) , .ZN( u1_u6_u5_n183 ) );
  INV_X1 u1_u6_u5_U29 (.A( u1_u6_u5_n123 ) , .ZN( u1_u6_u5_n185 ) );
  NOR2_X1 u1_u6_u5_U3 (.ZN( u1_u6_u5_n134 ) , .A1( u1_u6_u5_n183 ) , .A2( u1_u6_u5_n190 ) );
  INV_X1 u1_u6_u5_U30 (.A( u1_u6_u5_n161 ) , .ZN( u1_u6_u5_n184 ) );
  INV_X1 u1_u6_u5_U31 (.A( u1_u6_u5_n139 ) , .ZN( u1_u6_u5_n189 ) );
  INV_X1 u1_u6_u5_U32 (.A( u1_u6_u5_n157 ) , .ZN( u1_u6_u5_n190 ) );
  INV_X1 u1_u6_u5_U33 (.A( u1_u6_u5_n120 ) , .ZN( u1_u6_u5_n193 ) );
  NAND2_X1 u1_u6_u5_U34 (.ZN( u1_u6_u5_n111 ) , .A1( u1_u6_u5_n140 ) , .A2( u1_u6_u5_n155 ) );
  INV_X1 u1_u6_u5_U35 (.A( u1_u6_u5_n117 ) , .ZN( u1_u6_u5_n196 ) );
  OAI221_X1 u1_u6_u5_U36 (.A( u1_u6_u5_n116 ) , .ZN( u1_u6_u5_n117 ) , .B2( u1_u6_u5_n119 ) , .C1( u1_u6_u5_n153 ) , .C2( u1_u6_u5_n158 ) , .B1( u1_u6_u5_n172 ) );
  AOI222_X1 u1_u6_u5_U37 (.ZN( u1_u6_u5_n116 ) , .B2( u1_u6_u5_n145 ) , .C1( u1_u6_u5_n148 ) , .A2( u1_u6_u5_n174 ) , .C2( u1_u6_u5_n177 ) , .B1( u1_u6_u5_n187 ) , .A1( u1_u6_u5_n193 ) );
  INV_X1 u1_u6_u5_U38 (.A( u1_u6_u5_n115 ) , .ZN( u1_u6_u5_n187 ) );
  NOR2_X1 u1_u6_u5_U39 (.ZN( u1_u6_u5_n100 ) , .A1( u1_u6_u5_n170 ) , .A2( u1_u6_u5_n180 ) );
  INV_X1 u1_u6_u5_U4 (.A( u1_u6_u5_n138 ) , .ZN( u1_u6_u5_n191 ) );
  AOI22_X1 u1_u6_u5_U40 (.B2( u1_u6_u5_n131 ) , .A2( u1_u6_u5_n146 ) , .ZN( u1_u6_u5_n169 ) , .B1( u1_u6_u5_n174 ) , .A1( u1_u6_u5_n185 ) );
  NOR2_X1 u1_u6_u5_U41 (.A1( u1_u6_u5_n146 ) , .ZN( u1_u6_u5_n150 ) , .A2( u1_u6_u5_n173 ) );
  AOI21_X1 u1_u6_u5_U42 (.A( u1_u6_u5_n118 ) , .B2( u1_u6_u5_n145 ) , .ZN( u1_u6_u5_n168 ) , .B1( u1_u6_u5_n186 ) );
  INV_X1 u1_u6_u5_U43 (.A( u1_u6_u5_n122 ) , .ZN( u1_u6_u5_n186 ) );
  NOR2_X1 u1_u6_u5_U44 (.A1( u1_u6_u5_n146 ) , .ZN( u1_u6_u5_n152 ) , .A2( u1_u6_u5_n176 ) );
  NOR2_X1 u1_u6_u5_U45 (.A1( u1_u6_u5_n115 ) , .ZN( u1_u6_u5_n118 ) , .A2( u1_u6_u5_n153 ) );
  NOR2_X1 u1_u6_u5_U46 (.A2( u1_u6_u5_n145 ) , .ZN( u1_u6_u5_n156 ) , .A1( u1_u6_u5_n174 ) );
  NOR2_X1 u1_u6_u5_U47 (.ZN( u1_u6_u5_n121 ) , .A2( u1_u6_u5_n145 ) , .A1( u1_u6_u5_n176 ) );
  AOI22_X1 u1_u6_u5_U48 (.ZN( u1_u6_u5_n114 ) , .A2( u1_u6_u5_n137 ) , .A1( u1_u6_u5_n145 ) , .B2( u1_u6_u5_n175 ) , .B1( u1_u6_u5_n193 ) );
  OAI211_X1 u1_u6_u5_U49 (.B( u1_u6_u5_n124 ) , .A( u1_u6_u5_n125 ) , .C2( u1_u6_u5_n126 ) , .C1( u1_u6_u5_n127 ) , .ZN( u1_u6_u5_n128 ) );
  OAI21_X1 u1_u6_u5_U5 (.B2( u1_u6_u5_n136 ) , .B1( u1_u6_u5_n137 ) , .ZN( u1_u6_u5_n138 ) , .A( u1_u6_u5_n177 ) );
  NOR3_X1 u1_u6_u5_U50 (.ZN( u1_u6_u5_n127 ) , .A1( u1_u6_u5_n136 ) , .A3( u1_u6_u5_n148 ) , .A2( u1_u6_u5_n182 ) );
  OAI21_X1 u1_u6_u5_U51 (.ZN( u1_u6_u5_n124 ) , .A( u1_u6_u5_n177 ) , .B2( u1_u6_u5_n183 ) , .B1( u1_u6_u5_n189 ) );
  OAI21_X1 u1_u6_u5_U52 (.ZN( u1_u6_u5_n125 ) , .A( u1_u6_u5_n174 ) , .B2( u1_u6_u5_n185 ) , .B1( u1_u6_u5_n190 ) );
  AOI21_X1 u1_u6_u5_U53 (.A( u1_u6_u5_n153 ) , .B2( u1_u6_u5_n154 ) , .B1( u1_u6_u5_n155 ) , .ZN( u1_u6_u5_n164 ) );
  AOI21_X1 u1_u6_u5_U54 (.ZN( u1_u6_u5_n110 ) , .B1( u1_u6_u5_n122 ) , .B2( u1_u6_u5_n139 ) , .A( u1_u6_u5_n153 ) );
  INV_X1 u1_u6_u5_U55 (.A( u1_u6_u5_n153 ) , .ZN( u1_u6_u5_n176 ) );
  INV_X1 u1_u6_u5_U56 (.A( u1_u6_u5_n126 ) , .ZN( u1_u6_u5_n173 ) );
  AND2_X1 u1_u6_u5_U57 (.A2( u1_u6_u5_n104 ) , .A1( u1_u6_u5_n107 ) , .ZN( u1_u6_u5_n147 ) );
  AND2_X1 u1_u6_u5_U58 (.A2( u1_u6_u5_n104 ) , .A1( u1_u6_u5_n108 ) , .ZN( u1_u6_u5_n148 ) );
  NAND2_X1 u1_u6_u5_U59 (.A1( u1_u6_u5_n105 ) , .A2( u1_u6_u5_n106 ) , .ZN( u1_u6_u5_n158 ) );
  INV_X1 u1_u6_u5_U6 (.A( u1_u6_u5_n135 ) , .ZN( u1_u6_u5_n178 ) );
  NAND2_X1 u1_u6_u5_U60 (.A2( u1_u6_u5_n108 ) , .A1( u1_u6_u5_n109 ) , .ZN( u1_u6_u5_n139 ) );
  NAND2_X1 u1_u6_u5_U61 (.A1( u1_u6_u5_n106 ) , .A2( u1_u6_u5_n108 ) , .ZN( u1_u6_u5_n119 ) );
  NAND2_X1 u1_u6_u5_U62 (.A2( u1_u6_u5_n103 ) , .A1( u1_u6_u5_n105 ) , .ZN( u1_u6_u5_n140 ) );
  NAND2_X1 u1_u6_u5_U63 (.A2( u1_u6_u5_n104 ) , .A1( u1_u6_u5_n105 ) , .ZN( u1_u6_u5_n155 ) );
  NAND2_X1 u1_u6_u5_U64 (.A2( u1_u6_u5_n106 ) , .A1( u1_u6_u5_n107 ) , .ZN( u1_u6_u5_n122 ) );
  NAND2_X1 u1_u6_u5_U65 (.A2( u1_u6_u5_n100 ) , .A1( u1_u6_u5_n106 ) , .ZN( u1_u6_u5_n115 ) );
  NAND2_X1 u1_u6_u5_U66 (.A2( u1_u6_u5_n100 ) , .A1( u1_u6_u5_n103 ) , .ZN( u1_u6_u5_n161 ) );
  NAND2_X1 u1_u6_u5_U67 (.A1( u1_u6_u5_n105 ) , .A2( u1_u6_u5_n109 ) , .ZN( u1_u6_u5_n154 ) );
  INV_X1 u1_u6_u5_U68 (.A( u1_u6_u5_n146 ) , .ZN( u1_u6_u5_n172 ) );
  NAND2_X1 u1_u6_u5_U69 (.A1( u1_u6_u5_n103 ) , .A2( u1_u6_u5_n108 ) , .ZN( u1_u6_u5_n123 ) );
  OAI22_X1 u1_u6_u5_U7 (.B2( u1_u6_u5_n149 ) , .B1( u1_u6_u5_n150 ) , .A2( u1_u6_u5_n151 ) , .A1( u1_u6_u5_n152 ) , .ZN( u1_u6_u5_n165 ) );
  NAND2_X1 u1_u6_u5_U70 (.A2( u1_u6_u5_n103 ) , .A1( u1_u6_u5_n107 ) , .ZN( u1_u6_u5_n151 ) );
  NAND2_X1 u1_u6_u5_U71 (.A2( u1_u6_u5_n107 ) , .A1( u1_u6_u5_n109 ) , .ZN( u1_u6_u5_n120 ) );
  NAND2_X1 u1_u6_u5_U72 (.A2( u1_u6_u5_n100 ) , .A1( u1_u6_u5_n109 ) , .ZN( u1_u6_u5_n157 ) );
  AND2_X1 u1_u6_u5_U73 (.A2( u1_u6_u5_n100 ) , .A1( u1_u6_u5_n104 ) , .ZN( u1_u6_u5_n131 ) );
  INV_X1 u1_u6_u5_U74 (.A( u1_u6_u5_n102 ) , .ZN( u1_u6_u5_n195 ) );
  OAI221_X1 u1_u6_u5_U75 (.A( u1_u6_u5_n101 ) , .ZN( u1_u6_u5_n102 ) , .C2( u1_u6_u5_n115 ) , .C1( u1_u6_u5_n126 ) , .B1( u1_u6_u5_n134 ) , .B2( u1_u6_u5_n160 ) );
  OAI21_X1 u1_u6_u5_U76 (.ZN( u1_u6_u5_n101 ) , .B1( u1_u6_u5_n137 ) , .A( u1_u6_u5_n146 ) , .B2( u1_u6_u5_n147 ) );
  NOR2_X1 u1_u6_u5_U77 (.A2( u1_u6_X_34 ) , .A1( u1_u6_X_35 ) , .ZN( u1_u6_u5_n145 ) );
  NOR2_X1 u1_u6_u5_U78 (.A2( u1_u6_X_34 ) , .ZN( u1_u6_u5_n146 ) , .A1( u1_u6_u5_n171 ) );
  NOR2_X1 u1_u6_u5_U79 (.A2( u1_u6_X_31 ) , .A1( u1_u6_X_32 ) , .ZN( u1_u6_u5_n103 ) );
  NOR3_X1 u1_u6_u5_U8 (.A2( u1_u6_u5_n147 ) , .A1( u1_u6_u5_n148 ) , .ZN( u1_u6_u5_n149 ) , .A3( u1_u6_u5_n194 ) );
  NOR2_X1 u1_u6_u5_U80 (.A2( u1_u6_X_36 ) , .ZN( u1_u6_u5_n105 ) , .A1( u1_u6_u5_n180 ) );
  NOR2_X1 u1_u6_u5_U81 (.A2( u1_u6_X_33 ) , .ZN( u1_u6_u5_n108 ) , .A1( u1_u6_u5_n170 ) );
  NOR2_X1 u1_u6_u5_U82 (.A2( u1_u6_X_33 ) , .A1( u1_u6_X_36 ) , .ZN( u1_u6_u5_n107 ) );
  NOR2_X1 u1_u6_u5_U83 (.A2( u1_u6_X_31 ) , .ZN( u1_u6_u5_n104 ) , .A1( u1_u6_u5_n181 ) );
  NAND2_X1 u1_u6_u5_U84 (.A2( u1_u6_X_34 ) , .A1( u1_u6_X_35 ) , .ZN( u1_u6_u5_n153 ) );
  NAND2_X1 u1_u6_u5_U85 (.A1( u1_u6_X_34 ) , .ZN( u1_u6_u5_n126 ) , .A2( u1_u6_u5_n171 ) );
  AND2_X1 u1_u6_u5_U86 (.A1( u1_u6_X_31 ) , .A2( u1_u6_X_32 ) , .ZN( u1_u6_u5_n106 ) );
  AND2_X1 u1_u6_u5_U87 (.A1( u1_u6_X_31 ) , .ZN( u1_u6_u5_n109 ) , .A2( u1_u6_u5_n181 ) );
  INV_X1 u1_u6_u5_U88 (.A( u1_u6_X_33 ) , .ZN( u1_u6_u5_n180 ) );
  INV_X1 u1_u6_u5_U89 (.A( u1_u6_X_35 ) , .ZN( u1_u6_u5_n171 ) );
  NOR2_X1 u1_u6_u5_U9 (.ZN( u1_u6_u5_n135 ) , .A1( u1_u6_u5_n173 ) , .A2( u1_u6_u5_n176 ) );
  INV_X1 u1_u6_u5_U90 (.A( u1_u6_X_36 ) , .ZN( u1_u6_u5_n170 ) );
  INV_X1 u1_u6_u5_U91 (.A( u1_u6_X_32 ) , .ZN( u1_u6_u5_n181 ) );
  NAND4_X1 u1_u6_u5_U92 (.ZN( u1_out6_19 ) , .A4( u1_u6_u5_n166 ) , .A3( u1_u6_u5_n167 ) , .A2( u1_u6_u5_n168 ) , .A1( u1_u6_u5_n169 ) );
  AOI22_X1 u1_u6_u5_U93 (.B2( u1_u6_u5_n145 ) , .A2( u1_u6_u5_n146 ) , .ZN( u1_u6_u5_n167 ) , .B1( u1_u6_u5_n182 ) , .A1( u1_u6_u5_n189 ) );
  NOR4_X1 u1_u6_u5_U94 (.A4( u1_u6_u5_n162 ) , .A3( u1_u6_u5_n163 ) , .A2( u1_u6_u5_n164 ) , .A1( u1_u6_u5_n165 ) , .ZN( u1_u6_u5_n166 ) );
  NAND4_X1 u1_u6_u5_U95 (.ZN( u1_out6_29 ) , .A4( u1_u6_u5_n129 ) , .A3( u1_u6_u5_n130 ) , .A2( u1_u6_u5_n168 ) , .A1( u1_u6_u5_n196 ) );
  AOI221_X1 u1_u6_u5_U96 (.A( u1_u6_u5_n128 ) , .ZN( u1_u6_u5_n129 ) , .C2( u1_u6_u5_n132 ) , .B2( u1_u6_u5_n159 ) , .B1( u1_u6_u5_n176 ) , .C1( u1_u6_u5_n184 ) );
  AOI222_X1 u1_u6_u5_U97 (.ZN( u1_u6_u5_n130 ) , .A2( u1_u6_u5_n146 ) , .B1( u1_u6_u5_n147 ) , .C2( u1_u6_u5_n175 ) , .B2( u1_u6_u5_n179 ) , .A1( u1_u6_u5_n188 ) , .C1( u1_u6_u5_n194 ) );
  NAND4_X1 u1_u6_u5_U98 (.ZN( u1_out6_4 ) , .A4( u1_u6_u5_n112 ) , .A2( u1_u6_u5_n113 ) , .A1( u1_u6_u5_n114 ) , .A3( u1_u6_u5_n195 ) );
  AOI211_X1 u1_u6_u5_U99 (.A( u1_u6_u5_n110 ) , .C1( u1_u6_u5_n111 ) , .ZN( u1_u6_u5_n112 ) , .B( u1_u6_u5_n118 ) , .C2( u1_u6_u5_n177 ) );
  XOR2_X1 u1_u7_U20 (.B( u1_K8_36 ) , .A( u1_R6_25 ) , .Z( u1_u7_X_36 ) );
  XOR2_X1 u1_u7_U21 (.B( u1_K8_35 ) , .A( u1_R6_24 ) , .Z( u1_u7_X_35 ) );
  XOR2_X1 u1_u7_U22 (.B( u1_K8_34 ) , .A( u1_R6_23 ) , .Z( u1_u7_X_34 ) );
  XOR2_X1 u1_u7_U23 (.B( u1_K8_33 ) , .A( u1_R6_22 ) , .Z( u1_u7_X_33 ) );
  XOR2_X1 u1_u7_U24 (.B( u1_K8_32 ) , .A( u1_R6_21 ) , .Z( u1_u7_X_32 ) );
  XOR2_X1 u1_u7_U25 (.B( u1_K8_31 ) , .A( u1_R6_20 ) , .Z( u1_u7_X_31 ) );
  XOR2_X1 u1_u7_U26 (.B( u1_K8_30 ) , .A( u1_R6_21 ) , .Z( u1_u7_X_30 ) );
  XOR2_X1 u1_u7_U28 (.B( u1_K8_29 ) , .A( u1_R6_20 ) , .Z( u1_u7_X_29 ) );
  XOR2_X1 u1_u7_U29 (.B( u1_K8_28 ) , .A( u1_R6_19 ) , .Z( u1_u7_X_28 ) );
  XOR2_X1 u1_u7_U30 (.B( u1_K8_27 ) , .A( u1_R6_18 ) , .Z( u1_u7_X_27 ) );
  XOR2_X1 u1_u7_U31 (.B( u1_K8_26 ) , .A( u1_R6_17 ) , .Z( u1_u7_X_26 ) );
  XOR2_X1 u1_u7_U32 (.B( u1_K8_25 ) , .A( u1_R6_16 ) , .Z( u1_u7_X_25 ) );
  OAI22_X1 u1_u7_u4_U10 (.B2( u1_u7_u4_n135 ) , .ZN( u1_u7_u4_n137 ) , .B1( u1_u7_u4_n153 ) , .A1( u1_u7_u4_n155 ) , .A2( u1_u7_u4_n171 ) );
  AND3_X1 u1_u7_u4_U11 (.A2( u1_u7_u4_n134 ) , .ZN( u1_u7_u4_n135 ) , .A3( u1_u7_u4_n145 ) , .A1( u1_u7_u4_n157 ) );
  NAND2_X1 u1_u7_u4_U12 (.ZN( u1_u7_u4_n132 ) , .A2( u1_u7_u4_n170 ) , .A1( u1_u7_u4_n173 ) );
  AOI21_X1 u1_u7_u4_U13 (.B2( u1_u7_u4_n160 ) , .B1( u1_u7_u4_n161 ) , .ZN( u1_u7_u4_n162 ) , .A( u1_u7_u4_n170 ) );
  AOI21_X1 u1_u7_u4_U14 (.ZN( u1_u7_u4_n107 ) , .B2( u1_u7_u4_n143 ) , .A( u1_u7_u4_n174 ) , .B1( u1_u7_u4_n184 ) );
  AOI21_X1 u1_u7_u4_U15 (.B2( u1_u7_u4_n158 ) , .B1( u1_u7_u4_n159 ) , .ZN( u1_u7_u4_n163 ) , .A( u1_u7_u4_n174 ) );
  AOI21_X1 u1_u7_u4_U16 (.A( u1_u7_u4_n153 ) , .B2( u1_u7_u4_n154 ) , .B1( u1_u7_u4_n155 ) , .ZN( u1_u7_u4_n165 ) );
  AOI21_X1 u1_u7_u4_U17 (.A( u1_u7_u4_n156 ) , .B2( u1_u7_u4_n157 ) , .ZN( u1_u7_u4_n164 ) , .B1( u1_u7_u4_n184 ) );
  INV_X1 u1_u7_u4_U18 (.A( u1_u7_u4_n138 ) , .ZN( u1_u7_u4_n170 ) );
  AND2_X1 u1_u7_u4_U19 (.A2( u1_u7_u4_n120 ) , .ZN( u1_u7_u4_n155 ) , .A1( u1_u7_u4_n160 ) );
  INV_X1 u1_u7_u4_U20 (.A( u1_u7_u4_n156 ) , .ZN( u1_u7_u4_n175 ) );
  NAND2_X1 u1_u7_u4_U21 (.A2( u1_u7_u4_n118 ) , .ZN( u1_u7_u4_n131 ) , .A1( u1_u7_u4_n147 ) );
  NAND2_X1 u1_u7_u4_U22 (.A1( u1_u7_u4_n119 ) , .A2( u1_u7_u4_n120 ) , .ZN( u1_u7_u4_n130 ) );
  NAND2_X1 u1_u7_u4_U23 (.ZN( u1_u7_u4_n117 ) , .A2( u1_u7_u4_n118 ) , .A1( u1_u7_u4_n148 ) );
  NAND2_X1 u1_u7_u4_U24 (.ZN( u1_u7_u4_n129 ) , .A1( u1_u7_u4_n134 ) , .A2( u1_u7_u4_n148 ) );
  AND3_X1 u1_u7_u4_U25 (.A1( u1_u7_u4_n119 ) , .A2( u1_u7_u4_n143 ) , .A3( u1_u7_u4_n154 ) , .ZN( u1_u7_u4_n161 ) );
  AND2_X1 u1_u7_u4_U26 (.A1( u1_u7_u4_n145 ) , .A2( u1_u7_u4_n147 ) , .ZN( u1_u7_u4_n159 ) );
  OR3_X1 u1_u7_u4_U27 (.A3( u1_u7_u4_n114 ) , .A2( u1_u7_u4_n115 ) , .A1( u1_u7_u4_n116 ) , .ZN( u1_u7_u4_n136 ) );
  AOI21_X1 u1_u7_u4_U28 (.A( u1_u7_u4_n113 ) , .ZN( u1_u7_u4_n116 ) , .B2( u1_u7_u4_n173 ) , .B1( u1_u7_u4_n174 ) );
  AOI21_X1 u1_u7_u4_U29 (.ZN( u1_u7_u4_n115 ) , .B2( u1_u7_u4_n145 ) , .B1( u1_u7_u4_n146 ) , .A( u1_u7_u4_n156 ) );
  NOR2_X1 u1_u7_u4_U3 (.ZN( u1_u7_u4_n121 ) , .A1( u1_u7_u4_n181 ) , .A2( u1_u7_u4_n182 ) );
  OAI22_X1 u1_u7_u4_U30 (.ZN( u1_u7_u4_n114 ) , .A2( u1_u7_u4_n121 ) , .B1( u1_u7_u4_n160 ) , .B2( u1_u7_u4_n170 ) , .A1( u1_u7_u4_n171 ) );
  INV_X1 u1_u7_u4_U31 (.A( u1_u7_u4_n158 ) , .ZN( u1_u7_u4_n182 ) );
  INV_X1 u1_u7_u4_U32 (.ZN( u1_u7_u4_n181 ) , .A( u1_u7_u4_n96 ) );
  INV_X1 u1_u7_u4_U33 (.A( u1_u7_u4_n144 ) , .ZN( u1_u7_u4_n179 ) );
  INV_X1 u1_u7_u4_U34 (.A( u1_u7_u4_n157 ) , .ZN( u1_u7_u4_n178 ) );
  NAND2_X1 u1_u7_u4_U35 (.A2( u1_u7_u4_n154 ) , .A1( u1_u7_u4_n96 ) , .ZN( u1_u7_u4_n97 ) );
  INV_X1 u1_u7_u4_U36 (.ZN( u1_u7_u4_n186 ) , .A( u1_u7_u4_n95 ) );
  OAI221_X1 u1_u7_u4_U37 (.C1( u1_u7_u4_n134 ) , .B1( u1_u7_u4_n158 ) , .B2( u1_u7_u4_n171 ) , .C2( u1_u7_u4_n173 ) , .A( u1_u7_u4_n94 ) , .ZN( u1_u7_u4_n95 ) );
  AOI222_X1 u1_u7_u4_U38 (.B2( u1_u7_u4_n132 ) , .A1( u1_u7_u4_n138 ) , .C2( u1_u7_u4_n175 ) , .A2( u1_u7_u4_n179 ) , .C1( u1_u7_u4_n181 ) , .B1( u1_u7_u4_n185 ) , .ZN( u1_u7_u4_n94 ) );
  INV_X1 u1_u7_u4_U39 (.A( u1_u7_u4_n113 ) , .ZN( u1_u7_u4_n185 ) );
  INV_X1 u1_u7_u4_U4 (.A( u1_u7_u4_n117 ) , .ZN( u1_u7_u4_n184 ) );
  INV_X1 u1_u7_u4_U40 (.A( u1_u7_u4_n143 ) , .ZN( u1_u7_u4_n183 ) );
  NOR2_X1 u1_u7_u4_U41 (.ZN( u1_u7_u4_n138 ) , .A1( u1_u7_u4_n168 ) , .A2( u1_u7_u4_n169 ) );
  NOR2_X1 u1_u7_u4_U42 (.A1( u1_u7_u4_n150 ) , .A2( u1_u7_u4_n152 ) , .ZN( u1_u7_u4_n153 ) );
  NOR2_X1 u1_u7_u4_U43 (.A2( u1_u7_u4_n128 ) , .A1( u1_u7_u4_n138 ) , .ZN( u1_u7_u4_n156 ) );
  AOI22_X1 u1_u7_u4_U44 (.B2( u1_u7_u4_n122 ) , .A1( u1_u7_u4_n123 ) , .ZN( u1_u7_u4_n124 ) , .B1( u1_u7_u4_n128 ) , .A2( u1_u7_u4_n172 ) );
  NAND2_X1 u1_u7_u4_U45 (.A2( u1_u7_u4_n120 ) , .ZN( u1_u7_u4_n123 ) , .A1( u1_u7_u4_n161 ) );
  INV_X1 u1_u7_u4_U46 (.A( u1_u7_u4_n153 ) , .ZN( u1_u7_u4_n172 ) );
  AOI22_X1 u1_u7_u4_U47 (.B2( u1_u7_u4_n132 ) , .A2( u1_u7_u4_n133 ) , .ZN( u1_u7_u4_n140 ) , .A1( u1_u7_u4_n150 ) , .B1( u1_u7_u4_n179 ) );
  NAND2_X1 u1_u7_u4_U48 (.ZN( u1_u7_u4_n133 ) , .A2( u1_u7_u4_n146 ) , .A1( u1_u7_u4_n154 ) );
  NAND2_X1 u1_u7_u4_U49 (.A1( u1_u7_u4_n103 ) , .ZN( u1_u7_u4_n154 ) , .A2( u1_u7_u4_n98 ) );
  NOR4_X1 u1_u7_u4_U5 (.A4( u1_u7_u4_n106 ) , .A3( u1_u7_u4_n107 ) , .A2( u1_u7_u4_n108 ) , .A1( u1_u7_u4_n109 ) , .ZN( u1_u7_u4_n110 ) );
  NAND2_X1 u1_u7_u4_U50 (.A1( u1_u7_u4_n101 ) , .ZN( u1_u7_u4_n158 ) , .A2( u1_u7_u4_n99 ) );
  AOI21_X1 u1_u7_u4_U51 (.ZN( u1_u7_u4_n127 ) , .A( u1_u7_u4_n136 ) , .B2( u1_u7_u4_n150 ) , .B1( u1_u7_u4_n180 ) );
  INV_X1 u1_u7_u4_U52 (.A( u1_u7_u4_n160 ) , .ZN( u1_u7_u4_n180 ) );
  NAND2_X1 u1_u7_u4_U53 (.A2( u1_u7_u4_n104 ) , .A1( u1_u7_u4_n105 ) , .ZN( u1_u7_u4_n146 ) );
  NAND2_X1 u1_u7_u4_U54 (.A2( u1_u7_u4_n101 ) , .A1( u1_u7_u4_n102 ) , .ZN( u1_u7_u4_n160 ) );
  NAND2_X1 u1_u7_u4_U55 (.ZN( u1_u7_u4_n134 ) , .A1( u1_u7_u4_n98 ) , .A2( u1_u7_u4_n99 ) );
  NAND2_X1 u1_u7_u4_U56 (.A1( u1_u7_u4_n103 ) , .A2( u1_u7_u4_n104 ) , .ZN( u1_u7_u4_n143 ) );
  NAND2_X1 u1_u7_u4_U57 (.A2( u1_u7_u4_n105 ) , .ZN( u1_u7_u4_n145 ) , .A1( u1_u7_u4_n98 ) );
  NAND2_X1 u1_u7_u4_U58 (.A1( u1_u7_u4_n100 ) , .A2( u1_u7_u4_n105 ) , .ZN( u1_u7_u4_n120 ) );
  NAND2_X1 u1_u7_u4_U59 (.A1( u1_u7_u4_n102 ) , .A2( u1_u7_u4_n104 ) , .ZN( u1_u7_u4_n148 ) );
  AOI21_X1 u1_u7_u4_U6 (.ZN( u1_u7_u4_n106 ) , .B2( u1_u7_u4_n146 ) , .B1( u1_u7_u4_n158 ) , .A( u1_u7_u4_n170 ) );
  NAND2_X1 u1_u7_u4_U60 (.A2( u1_u7_u4_n100 ) , .A1( u1_u7_u4_n103 ) , .ZN( u1_u7_u4_n157 ) );
  INV_X1 u1_u7_u4_U61 (.A( u1_u7_u4_n150 ) , .ZN( u1_u7_u4_n173 ) );
  INV_X1 u1_u7_u4_U62 (.A( u1_u7_u4_n152 ) , .ZN( u1_u7_u4_n171 ) );
  NAND2_X1 u1_u7_u4_U63 (.A1( u1_u7_u4_n100 ) , .ZN( u1_u7_u4_n118 ) , .A2( u1_u7_u4_n99 ) );
  NAND2_X1 u1_u7_u4_U64 (.A2( u1_u7_u4_n100 ) , .A1( u1_u7_u4_n102 ) , .ZN( u1_u7_u4_n144 ) );
  NAND2_X1 u1_u7_u4_U65 (.A2( u1_u7_u4_n101 ) , .A1( u1_u7_u4_n105 ) , .ZN( u1_u7_u4_n96 ) );
  INV_X1 u1_u7_u4_U66 (.A( u1_u7_u4_n128 ) , .ZN( u1_u7_u4_n174 ) );
  NAND2_X1 u1_u7_u4_U67 (.A2( u1_u7_u4_n102 ) , .ZN( u1_u7_u4_n119 ) , .A1( u1_u7_u4_n98 ) );
  NAND2_X1 u1_u7_u4_U68 (.A2( u1_u7_u4_n101 ) , .A1( u1_u7_u4_n103 ) , .ZN( u1_u7_u4_n147 ) );
  NAND2_X1 u1_u7_u4_U69 (.A2( u1_u7_u4_n104 ) , .ZN( u1_u7_u4_n113 ) , .A1( u1_u7_u4_n99 ) );
  AOI21_X1 u1_u7_u4_U7 (.ZN( u1_u7_u4_n108 ) , .B2( u1_u7_u4_n134 ) , .B1( u1_u7_u4_n155 ) , .A( u1_u7_u4_n156 ) );
  NOR2_X1 u1_u7_u4_U70 (.A2( u1_u7_X_28 ) , .ZN( u1_u7_u4_n150 ) , .A1( u1_u7_u4_n168 ) );
  NOR2_X1 u1_u7_u4_U71 (.A2( u1_u7_X_29 ) , .ZN( u1_u7_u4_n152 ) , .A1( u1_u7_u4_n169 ) );
  NOR2_X1 u1_u7_u4_U72 (.A2( u1_u7_X_26 ) , .ZN( u1_u7_u4_n100 ) , .A1( u1_u7_u4_n177 ) );
  NOR2_X1 u1_u7_u4_U73 (.A2( u1_u7_X_30 ) , .ZN( u1_u7_u4_n105 ) , .A1( u1_u7_u4_n176 ) );
  NOR2_X1 u1_u7_u4_U74 (.A2( u1_u7_X_28 ) , .A1( u1_u7_X_29 ) , .ZN( u1_u7_u4_n128 ) );
  NOR2_X1 u1_u7_u4_U75 (.A2( u1_u7_X_25 ) , .A1( u1_u7_X_26 ) , .ZN( u1_u7_u4_n98 ) );
  NOR2_X1 u1_u7_u4_U76 (.A2( u1_u7_X_27 ) , .A1( u1_u7_X_30 ) , .ZN( u1_u7_u4_n102 ) );
  AND2_X1 u1_u7_u4_U77 (.A2( u1_u7_X_25 ) , .A1( u1_u7_X_26 ) , .ZN( u1_u7_u4_n104 ) );
  AND2_X1 u1_u7_u4_U78 (.A1( u1_u7_X_30 ) , .A2( u1_u7_u4_n176 ) , .ZN( u1_u7_u4_n99 ) );
  AND2_X1 u1_u7_u4_U79 (.A1( u1_u7_X_26 ) , .ZN( u1_u7_u4_n101 ) , .A2( u1_u7_u4_n177 ) );
  AOI21_X1 u1_u7_u4_U8 (.ZN( u1_u7_u4_n109 ) , .A( u1_u7_u4_n153 ) , .B1( u1_u7_u4_n159 ) , .B2( u1_u7_u4_n184 ) );
  AND2_X1 u1_u7_u4_U80 (.A1( u1_u7_X_27 ) , .A2( u1_u7_X_30 ) , .ZN( u1_u7_u4_n103 ) );
  INV_X1 u1_u7_u4_U81 (.A( u1_u7_X_28 ) , .ZN( u1_u7_u4_n169 ) );
  INV_X1 u1_u7_u4_U82 (.A( u1_u7_X_29 ) , .ZN( u1_u7_u4_n168 ) );
  INV_X1 u1_u7_u4_U83 (.A( u1_u7_X_25 ) , .ZN( u1_u7_u4_n177 ) );
  INV_X1 u1_u7_u4_U84 (.A( u1_u7_X_27 ) , .ZN( u1_u7_u4_n176 ) );
  NAND4_X1 u1_u7_u4_U85 (.ZN( u1_out7_25 ) , .A4( u1_u7_u4_n139 ) , .A3( u1_u7_u4_n140 ) , .A2( u1_u7_u4_n141 ) , .A1( u1_u7_u4_n142 ) );
  OAI21_X1 u1_u7_u4_U86 (.A( u1_u7_u4_n128 ) , .B2( u1_u7_u4_n129 ) , .B1( u1_u7_u4_n130 ) , .ZN( u1_u7_u4_n142 ) );
  OAI21_X1 u1_u7_u4_U87 (.B2( u1_u7_u4_n131 ) , .ZN( u1_u7_u4_n141 ) , .A( u1_u7_u4_n175 ) , .B1( u1_u7_u4_n183 ) );
  NAND4_X1 u1_u7_u4_U88 (.ZN( u1_out7_14 ) , .A4( u1_u7_u4_n124 ) , .A3( u1_u7_u4_n125 ) , .A2( u1_u7_u4_n126 ) , .A1( u1_u7_u4_n127 ) );
  AOI22_X1 u1_u7_u4_U89 (.B2( u1_u7_u4_n117 ) , .ZN( u1_u7_u4_n126 ) , .A1( u1_u7_u4_n129 ) , .B1( u1_u7_u4_n152 ) , .A2( u1_u7_u4_n175 ) );
  AOI211_X1 u1_u7_u4_U9 (.B( u1_u7_u4_n136 ) , .A( u1_u7_u4_n137 ) , .C2( u1_u7_u4_n138 ) , .ZN( u1_u7_u4_n139 ) , .C1( u1_u7_u4_n182 ) );
  AOI22_X1 u1_u7_u4_U90 (.ZN( u1_u7_u4_n125 ) , .B2( u1_u7_u4_n131 ) , .A2( u1_u7_u4_n132 ) , .B1( u1_u7_u4_n138 ) , .A1( u1_u7_u4_n178 ) );
  NAND4_X1 u1_u7_u4_U91 (.ZN( u1_out7_8 ) , .A4( u1_u7_u4_n110 ) , .A3( u1_u7_u4_n111 ) , .A2( u1_u7_u4_n112 ) , .A1( u1_u7_u4_n186 ) );
  NAND2_X1 u1_u7_u4_U92 (.ZN( u1_u7_u4_n112 ) , .A2( u1_u7_u4_n130 ) , .A1( u1_u7_u4_n150 ) );
  AOI22_X1 u1_u7_u4_U93 (.ZN( u1_u7_u4_n111 ) , .B2( u1_u7_u4_n132 ) , .A1( u1_u7_u4_n152 ) , .B1( u1_u7_u4_n178 ) , .A2( u1_u7_u4_n97 ) );
  AOI22_X1 u1_u7_u4_U94 (.B2( u1_u7_u4_n149 ) , .B1( u1_u7_u4_n150 ) , .A2( u1_u7_u4_n151 ) , .A1( u1_u7_u4_n152 ) , .ZN( u1_u7_u4_n167 ) );
  NOR4_X1 u1_u7_u4_U95 (.A4( u1_u7_u4_n162 ) , .A3( u1_u7_u4_n163 ) , .A2( u1_u7_u4_n164 ) , .A1( u1_u7_u4_n165 ) , .ZN( u1_u7_u4_n166 ) );
  NAND3_X1 u1_u7_u4_U96 (.ZN( u1_out7_3 ) , .A3( u1_u7_u4_n166 ) , .A1( u1_u7_u4_n167 ) , .A2( u1_u7_u4_n186 ) );
  NAND3_X1 u1_u7_u4_U97 (.A3( u1_u7_u4_n146 ) , .A2( u1_u7_u4_n147 ) , .A1( u1_u7_u4_n148 ) , .ZN( u1_u7_u4_n149 ) );
  NAND3_X1 u1_u7_u4_U98 (.A3( u1_u7_u4_n143 ) , .A2( u1_u7_u4_n144 ) , .A1( u1_u7_u4_n145 ) , .ZN( u1_u7_u4_n151 ) );
  NAND3_X1 u1_u7_u4_U99 (.A3( u1_u7_u4_n121 ) , .ZN( u1_u7_u4_n122 ) , .A2( u1_u7_u4_n144 ) , .A1( u1_u7_u4_n154 ) );
  INV_X1 u1_u7_u5_U10 (.A( u1_u7_u5_n121 ) , .ZN( u1_u7_u5_n177 ) );
  NOR3_X1 u1_u7_u5_U100 (.A3( u1_u7_u5_n141 ) , .A1( u1_u7_u5_n142 ) , .ZN( u1_u7_u5_n143 ) , .A2( u1_u7_u5_n191 ) );
  NAND4_X1 u1_u7_u5_U101 (.ZN( u1_out7_4 ) , .A4( u1_u7_u5_n112 ) , .A2( u1_u7_u5_n113 ) , .A1( u1_u7_u5_n114 ) , .A3( u1_u7_u5_n195 ) );
  AOI211_X1 u1_u7_u5_U102 (.A( u1_u7_u5_n110 ) , .C1( u1_u7_u5_n111 ) , .ZN( u1_u7_u5_n112 ) , .B( u1_u7_u5_n118 ) , .C2( u1_u7_u5_n177 ) );
  AOI222_X1 u1_u7_u5_U103 (.ZN( u1_u7_u5_n113 ) , .A1( u1_u7_u5_n131 ) , .C1( u1_u7_u5_n148 ) , .B2( u1_u7_u5_n174 ) , .C2( u1_u7_u5_n178 ) , .A2( u1_u7_u5_n179 ) , .B1( u1_u7_u5_n99 ) );
  NAND3_X1 u1_u7_u5_U104 (.A2( u1_u7_u5_n154 ) , .A3( u1_u7_u5_n158 ) , .A1( u1_u7_u5_n161 ) , .ZN( u1_u7_u5_n99 ) );
  NOR2_X1 u1_u7_u5_U11 (.ZN( u1_u7_u5_n160 ) , .A2( u1_u7_u5_n173 ) , .A1( u1_u7_u5_n177 ) );
  INV_X1 u1_u7_u5_U12 (.A( u1_u7_u5_n150 ) , .ZN( u1_u7_u5_n174 ) );
  AOI21_X1 u1_u7_u5_U13 (.A( u1_u7_u5_n160 ) , .B2( u1_u7_u5_n161 ) , .ZN( u1_u7_u5_n162 ) , .B1( u1_u7_u5_n192 ) );
  INV_X1 u1_u7_u5_U14 (.A( u1_u7_u5_n159 ) , .ZN( u1_u7_u5_n192 ) );
  AOI21_X1 u1_u7_u5_U15 (.A( u1_u7_u5_n156 ) , .B2( u1_u7_u5_n157 ) , .B1( u1_u7_u5_n158 ) , .ZN( u1_u7_u5_n163 ) );
  AOI21_X1 u1_u7_u5_U16 (.B2( u1_u7_u5_n139 ) , .B1( u1_u7_u5_n140 ) , .ZN( u1_u7_u5_n141 ) , .A( u1_u7_u5_n150 ) );
  OAI21_X1 u1_u7_u5_U17 (.A( u1_u7_u5_n133 ) , .B2( u1_u7_u5_n134 ) , .B1( u1_u7_u5_n135 ) , .ZN( u1_u7_u5_n142 ) );
  OAI21_X1 u1_u7_u5_U18 (.ZN( u1_u7_u5_n133 ) , .B2( u1_u7_u5_n147 ) , .A( u1_u7_u5_n173 ) , .B1( u1_u7_u5_n188 ) );
  NAND2_X1 u1_u7_u5_U19 (.A2( u1_u7_u5_n119 ) , .A1( u1_u7_u5_n123 ) , .ZN( u1_u7_u5_n137 ) );
  INV_X1 u1_u7_u5_U20 (.A( u1_u7_u5_n155 ) , .ZN( u1_u7_u5_n194 ) );
  NAND2_X1 u1_u7_u5_U21 (.A1( u1_u7_u5_n121 ) , .ZN( u1_u7_u5_n132 ) , .A2( u1_u7_u5_n172 ) );
  NAND2_X1 u1_u7_u5_U22 (.A2( u1_u7_u5_n122 ) , .ZN( u1_u7_u5_n136 ) , .A1( u1_u7_u5_n154 ) );
  NAND2_X1 u1_u7_u5_U23 (.A2( u1_u7_u5_n119 ) , .A1( u1_u7_u5_n120 ) , .ZN( u1_u7_u5_n159 ) );
  INV_X1 u1_u7_u5_U24 (.A( u1_u7_u5_n156 ) , .ZN( u1_u7_u5_n175 ) );
  INV_X1 u1_u7_u5_U25 (.A( u1_u7_u5_n158 ) , .ZN( u1_u7_u5_n188 ) );
  INV_X1 u1_u7_u5_U26 (.A( u1_u7_u5_n152 ) , .ZN( u1_u7_u5_n179 ) );
  INV_X1 u1_u7_u5_U27 (.A( u1_u7_u5_n140 ) , .ZN( u1_u7_u5_n182 ) );
  INV_X1 u1_u7_u5_U28 (.A( u1_u7_u5_n151 ) , .ZN( u1_u7_u5_n183 ) );
  INV_X1 u1_u7_u5_U29 (.A( u1_u7_u5_n123 ) , .ZN( u1_u7_u5_n185 ) );
  NOR2_X1 u1_u7_u5_U3 (.ZN( u1_u7_u5_n134 ) , .A1( u1_u7_u5_n183 ) , .A2( u1_u7_u5_n190 ) );
  INV_X1 u1_u7_u5_U30 (.A( u1_u7_u5_n161 ) , .ZN( u1_u7_u5_n184 ) );
  INV_X1 u1_u7_u5_U31 (.A( u1_u7_u5_n139 ) , .ZN( u1_u7_u5_n189 ) );
  INV_X1 u1_u7_u5_U32 (.A( u1_u7_u5_n157 ) , .ZN( u1_u7_u5_n190 ) );
  INV_X1 u1_u7_u5_U33 (.A( u1_u7_u5_n120 ) , .ZN( u1_u7_u5_n193 ) );
  NAND2_X1 u1_u7_u5_U34 (.ZN( u1_u7_u5_n111 ) , .A1( u1_u7_u5_n140 ) , .A2( u1_u7_u5_n155 ) );
  NOR2_X1 u1_u7_u5_U35 (.ZN( u1_u7_u5_n100 ) , .A1( u1_u7_u5_n170 ) , .A2( u1_u7_u5_n180 ) );
  INV_X1 u1_u7_u5_U36 (.A( u1_u7_u5_n117 ) , .ZN( u1_u7_u5_n196 ) );
  OAI221_X1 u1_u7_u5_U37 (.A( u1_u7_u5_n116 ) , .ZN( u1_u7_u5_n117 ) , .B2( u1_u7_u5_n119 ) , .C1( u1_u7_u5_n153 ) , .C2( u1_u7_u5_n158 ) , .B1( u1_u7_u5_n172 ) );
  AOI222_X1 u1_u7_u5_U38 (.ZN( u1_u7_u5_n116 ) , .B2( u1_u7_u5_n145 ) , .C1( u1_u7_u5_n148 ) , .A2( u1_u7_u5_n174 ) , .C2( u1_u7_u5_n177 ) , .B1( u1_u7_u5_n187 ) , .A1( u1_u7_u5_n193 ) );
  INV_X1 u1_u7_u5_U39 (.A( u1_u7_u5_n115 ) , .ZN( u1_u7_u5_n187 ) );
  INV_X1 u1_u7_u5_U4 (.A( u1_u7_u5_n138 ) , .ZN( u1_u7_u5_n191 ) );
  AOI22_X1 u1_u7_u5_U40 (.B2( u1_u7_u5_n131 ) , .A2( u1_u7_u5_n146 ) , .ZN( u1_u7_u5_n169 ) , .B1( u1_u7_u5_n174 ) , .A1( u1_u7_u5_n185 ) );
  NOR2_X1 u1_u7_u5_U41 (.A1( u1_u7_u5_n146 ) , .ZN( u1_u7_u5_n150 ) , .A2( u1_u7_u5_n173 ) );
  AOI21_X1 u1_u7_u5_U42 (.A( u1_u7_u5_n118 ) , .B2( u1_u7_u5_n145 ) , .ZN( u1_u7_u5_n168 ) , .B1( u1_u7_u5_n186 ) );
  INV_X1 u1_u7_u5_U43 (.A( u1_u7_u5_n122 ) , .ZN( u1_u7_u5_n186 ) );
  NOR2_X1 u1_u7_u5_U44 (.A1( u1_u7_u5_n146 ) , .ZN( u1_u7_u5_n152 ) , .A2( u1_u7_u5_n176 ) );
  NOR2_X1 u1_u7_u5_U45 (.A1( u1_u7_u5_n115 ) , .ZN( u1_u7_u5_n118 ) , .A2( u1_u7_u5_n153 ) );
  NOR2_X1 u1_u7_u5_U46 (.A2( u1_u7_u5_n145 ) , .ZN( u1_u7_u5_n156 ) , .A1( u1_u7_u5_n174 ) );
  NOR2_X1 u1_u7_u5_U47 (.ZN( u1_u7_u5_n121 ) , .A2( u1_u7_u5_n145 ) , .A1( u1_u7_u5_n176 ) );
  AOI22_X1 u1_u7_u5_U48 (.ZN( u1_u7_u5_n114 ) , .A2( u1_u7_u5_n137 ) , .A1( u1_u7_u5_n145 ) , .B2( u1_u7_u5_n175 ) , .B1( u1_u7_u5_n193 ) );
  OAI211_X1 u1_u7_u5_U49 (.B( u1_u7_u5_n124 ) , .A( u1_u7_u5_n125 ) , .C2( u1_u7_u5_n126 ) , .C1( u1_u7_u5_n127 ) , .ZN( u1_u7_u5_n128 ) );
  OAI21_X1 u1_u7_u5_U5 (.B2( u1_u7_u5_n136 ) , .B1( u1_u7_u5_n137 ) , .ZN( u1_u7_u5_n138 ) , .A( u1_u7_u5_n177 ) );
  NOR3_X1 u1_u7_u5_U50 (.ZN( u1_u7_u5_n127 ) , .A1( u1_u7_u5_n136 ) , .A3( u1_u7_u5_n148 ) , .A2( u1_u7_u5_n182 ) );
  OAI21_X1 u1_u7_u5_U51 (.ZN( u1_u7_u5_n124 ) , .A( u1_u7_u5_n177 ) , .B2( u1_u7_u5_n183 ) , .B1( u1_u7_u5_n189 ) );
  OAI21_X1 u1_u7_u5_U52 (.ZN( u1_u7_u5_n125 ) , .A( u1_u7_u5_n174 ) , .B2( u1_u7_u5_n185 ) , .B1( u1_u7_u5_n190 ) );
  AOI21_X1 u1_u7_u5_U53 (.A( u1_u7_u5_n153 ) , .B2( u1_u7_u5_n154 ) , .B1( u1_u7_u5_n155 ) , .ZN( u1_u7_u5_n164 ) );
  AOI21_X1 u1_u7_u5_U54 (.ZN( u1_u7_u5_n110 ) , .B1( u1_u7_u5_n122 ) , .B2( u1_u7_u5_n139 ) , .A( u1_u7_u5_n153 ) );
  INV_X1 u1_u7_u5_U55 (.A( u1_u7_u5_n153 ) , .ZN( u1_u7_u5_n176 ) );
  INV_X1 u1_u7_u5_U56 (.A( u1_u7_u5_n126 ) , .ZN( u1_u7_u5_n173 ) );
  AND2_X1 u1_u7_u5_U57 (.A2( u1_u7_u5_n104 ) , .A1( u1_u7_u5_n107 ) , .ZN( u1_u7_u5_n147 ) );
  AND2_X1 u1_u7_u5_U58 (.A2( u1_u7_u5_n104 ) , .A1( u1_u7_u5_n108 ) , .ZN( u1_u7_u5_n148 ) );
  NAND2_X1 u1_u7_u5_U59 (.A1( u1_u7_u5_n105 ) , .A2( u1_u7_u5_n106 ) , .ZN( u1_u7_u5_n158 ) );
  INV_X1 u1_u7_u5_U6 (.A( u1_u7_u5_n135 ) , .ZN( u1_u7_u5_n178 ) );
  NAND2_X1 u1_u7_u5_U60 (.A2( u1_u7_u5_n108 ) , .A1( u1_u7_u5_n109 ) , .ZN( u1_u7_u5_n139 ) );
  NAND2_X1 u1_u7_u5_U61 (.A1( u1_u7_u5_n106 ) , .A2( u1_u7_u5_n108 ) , .ZN( u1_u7_u5_n119 ) );
  NAND2_X1 u1_u7_u5_U62 (.A2( u1_u7_u5_n103 ) , .A1( u1_u7_u5_n105 ) , .ZN( u1_u7_u5_n140 ) );
  NAND2_X1 u1_u7_u5_U63 (.A2( u1_u7_u5_n104 ) , .A1( u1_u7_u5_n105 ) , .ZN( u1_u7_u5_n155 ) );
  NAND2_X1 u1_u7_u5_U64 (.A2( u1_u7_u5_n106 ) , .A1( u1_u7_u5_n107 ) , .ZN( u1_u7_u5_n122 ) );
  NAND2_X1 u1_u7_u5_U65 (.A2( u1_u7_u5_n100 ) , .A1( u1_u7_u5_n106 ) , .ZN( u1_u7_u5_n115 ) );
  NAND2_X1 u1_u7_u5_U66 (.A2( u1_u7_u5_n100 ) , .A1( u1_u7_u5_n103 ) , .ZN( u1_u7_u5_n161 ) );
  NAND2_X1 u1_u7_u5_U67 (.A1( u1_u7_u5_n105 ) , .A2( u1_u7_u5_n109 ) , .ZN( u1_u7_u5_n154 ) );
  INV_X1 u1_u7_u5_U68 (.A( u1_u7_u5_n146 ) , .ZN( u1_u7_u5_n172 ) );
  NAND2_X1 u1_u7_u5_U69 (.A1( u1_u7_u5_n103 ) , .A2( u1_u7_u5_n108 ) , .ZN( u1_u7_u5_n123 ) );
  OAI22_X1 u1_u7_u5_U7 (.B2( u1_u7_u5_n149 ) , .B1( u1_u7_u5_n150 ) , .A2( u1_u7_u5_n151 ) , .A1( u1_u7_u5_n152 ) , .ZN( u1_u7_u5_n165 ) );
  NAND2_X1 u1_u7_u5_U70 (.A2( u1_u7_u5_n103 ) , .A1( u1_u7_u5_n107 ) , .ZN( u1_u7_u5_n151 ) );
  NAND2_X1 u1_u7_u5_U71 (.A2( u1_u7_u5_n107 ) , .A1( u1_u7_u5_n109 ) , .ZN( u1_u7_u5_n120 ) );
  NAND2_X1 u1_u7_u5_U72 (.A2( u1_u7_u5_n100 ) , .A1( u1_u7_u5_n109 ) , .ZN( u1_u7_u5_n157 ) );
  AND2_X1 u1_u7_u5_U73 (.A2( u1_u7_u5_n100 ) , .A1( u1_u7_u5_n104 ) , .ZN( u1_u7_u5_n131 ) );
  INV_X1 u1_u7_u5_U74 (.A( u1_u7_u5_n102 ) , .ZN( u1_u7_u5_n195 ) );
  OAI221_X1 u1_u7_u5_U75 (.A( u1_u7_u5_n101 ) , .ZN( u1_u7_u5_n102 ) , .C2( u1_u7_u5_n115 ) , .C1( u1_u7_u5_n126 ) , .B1( u1_u7_u5_n134 ) , .B2( u1_u7_u5_n160 ) );
  OAI21_X1 u1_u7_u5_U76 (.ZN( u1_u7_u5_n101 ) , .B1( u1_u7_u5_n137 ) , .A( u1_u7_u5_n146 ) , .B2( u1_u7_u5_n147 ) );
  NOR2_X1 u1_u7_u5_U77 (.A2( u1_u7_X_34 ) , .A1( u1_u7_X_35 ) , .ZN( u1_u7_u5_n145 ) );
  NOR2_X1 u1_u7_u5_U78 (.A2( u1_u7_X_34 ) , .ZN( u1_u7_u5_n146 ) , .A1( u1_u7_u5_n171 ) );
  NOR2_X1 u1_u7_u5_U79 (.A2( u1_u7_X_31 ) , .A1( u1_u7_X_32 ) , .ZN( u1_u7_u5_n103 ) );
  NOR3_X1 u1_u7_u5_U8 (.A2( u1_u7_u5_n147 ) , .A1( u1_u7_u5_n148 ) , .ZN( u1_u7_u5_n149 ) , .A3( u1_u7_u5_n194 ) );
  NOR2_X1 u1_u7_u5_U80 (.A2( u1_u7_X_36 ) , .ZN( u1_u7_u5_n105 ) , .A1( u1_u7_u5_n180 ) );
  NOR2_X1 u1_u7_u5_U81 (.A2( u1_u7_X_33 ) , .ZN( u1_u7_u5_n108 ) , .A1( u1_u7_u5_n170 ) );
  NOR2_X1 u1_u7_u5_U82 (.A2( u1_u7_X_33 ) , .A1( u1_u7_X_36 ) , .ZN( u1_u7_u5_n107 ) );
  NOR2_X1 u1_u7_u5_U83 (.A2( u1_u7_X_31 ) , .ZN( u1_u7_u5_n104 ) , .A1( u1_u7_u5_n181 ) );
  NAND2_X1 u1_u7_u5_U84 (.A2( u1_u7_X_34 ) , .A1( u1_u7_X_35 ) , .ZN( u1_u7_u5_n153 ) );
  NAND2_X1 u1_u7_u5_U85 (.A1( u1_u7_X_34 ) , .ZN( u1_u7_u5_n126 ) , .A2( u1_u7_u5_n171 ) );
  AND2_X1 u1_u7_u5_U86 (.A1( u1_u7_X_31 ) , .A2( u1_u7_X_32 ) , .ZN( u1_u7_u5_n106 ) );
  AND2_X1 u1_u7_u5_U87 (.A1( u1_u7_X_31 ) , .ZN( u1_u7_u5_n109 ) , .A2( u1_u7_u5_n181 ) );
  INV_X1 u1_u7_u5_U88 (.A( u1_u7_X_33 ) , .ZN( u1_u7_u5_n180 ) );
  INV_X1 u1_u7_u5_U89 (.A( u1_u7_X_35 ) , .ZN( u1_u7_u5_n171 ) );
  NOR2_X1 u1_u7_u5_U9 (.ZN( u1_u7_u5_n135 ) , .A1( u1_u7_u5_n173 ) , .A2( u1_u7_u5_n176 ) );
  INV_X1 u1_u7_u5_U90 (.A( u1_u7_X_36 ) , .ZN( u1_u7_u5_n170 ) );
  INV_X1 u1_u7_u5_U91 (.A( u1_u7_X_32 ) , .ZN( u1_u7_u5_n181 ) );
  NAND4_X1 u1_u7_u5_U92 (.ZN( u1_out7_29 ) , .A4( u1_u7_u5_n129 ) , .A3( u1_u7_u5_n130 ) , .A2( u1_u7_u5_n168 ) , .A1( u1_u7_u5_n196 ) );
  AOI221_X1 u1_u7_u5_U93 (.A( u1_u7_u5_n128 ) , .ZN( u1_u7_u5_n129 ) , .C2( u1_u7_u5_n132 ) , .B2( u1_u7_u5_n159 ) , .B1( u1_u7_u5_n176 ) , .C1( u1_u7_u5_n184 ) );
  AOI222_X1 u1_u7_u5_U94 (.ZN( u1_u7_u5_n130 ) , .A2( u1_u7_u5_n146 ) , .B1( u1_u7_u5_n147 ) , .C2( u1_u7_u5_n175 ) , .B2( u1_u7_u5_n179 ) , .A1( u1_u7_u5_n188 ) , .C1( u1_u7_u5_n194 ) );
  NAND4_X1 u1_u7_u5_U95 (.ZN( u1_out7_19 ) , .A4( u1_u7_u5_n166 ) , .A3( u1_u7_u5_n167 ) , .A2( u1_u7_u5_n168 ) , .A1( u1_u7_u5_n169 ) );
  AOI22_X1 u1_u7_u5_U96 (.B2( u1_u7_u5_n145 ) , .A2( u1_u7_u5_n146 ) , .ZN( u1_u7_u5_n167 ) , .B1( u1_u7_u5_n182 ) , .A1( u1_u7_u5_n189 ) );
  NOR4_X1 u1_u7_u5_U97 (.A4( u1_u7_u5_n162 ) , .A3( u1_u7_u5_n163 ) , .A2( u1_u7_u5_n164 ) , .A1( u1_u7_u5_n165 ) , .ZN( u1_u7_u5_n166 ) );
  NAND4_X1 u1_u7_u5_U98 (.ZN( u1_out7_11 ) , .A4( u1_u7_u5_n143 ) , .A3( u1_u7_u5_n144 ) , .A2( u1_u7_u5_n169 ) , .A1( u1_u7_u5_n196 ) );
  AOI22_X1 u1_u7_u5_U99 (.A2( u1_u7_u5_n132 ) , .ZN( u1_u7_u5_n144 ) , .B2( u1_u7_u5_n145 ) , .B1( u1_u7_u5_n184 ) , .A1( u1_u7_u5_n194 ) );
  XOR2_X1 u1_u8_U26 (.B( u1_K9_30 ) , .A( u1_R7_21 ) , .Z( u1_u8_X_30 ) );
  XOR2_X1 u1_u8_U28 (.B( u1_K9_29 ) , .A( u1_R7_20 ) , .Z( u1_u8_X_29 ) );
  XOR2_X1 u1_u8_U29 (.B( u1_K9_28 ) , .A( u1_R7_19 ) , .Z( u1_u8_X_28 ) );
  XOR2_X1 u1_u8_U30 (.B( u1_K9_27 ) , .A( u1_R7_18 ) , .Z( u1_u8_X_27 ) );
  XOR2_X1 u1_u8_U31 (.B( u1_K9_26 ) , .A( u1_R7_17 ) , .Z( u1_u8_X_26 ) );
  XOR2_X1 u1_u8_U32 (.B( u1_K9_25 ) , .A( u1_R7_16 ) , .Z( u1_u8_X_25 ) );
  OAI22_X1 u1_u8_u4_U10 (.B2( u1_u8_u4_n135 ) , .ZN( u1_u8_u4_n137 ) , .B1( u1_u8_u4_n153 ) , .A1( u1_u8_u4_n155 ) , .A2( u1_u8_u4_n171 ) );
  AND3_X1 u1_u8_u4_U11 (.A2( u1_u8_u4_n134 ) , .ZN( u1_u8_u4_n135 ) , .A3( u1_u8_u4_n145 ) , .A1( u1_u8_u4_n157 ) );
  NAND2_X1 u1_u8_u4_U12 (.ZN( u1_u8_u4_n132 ) , .A2( u1_u8_u4_n170 ) , .A1( u1_u8_u4_n173 ) );
  AOI21_X1 u1_u8_u4_U13 (.B2( u1_u8_u4_n160 ) , .B1( u1_u8_u4_n161 ) , .ZN( u1_u8_u4_n162 ) , .A( u1_u8_u4_n170 ) );
  AOI21_X1 u1_u8_u4_U14 (.ZN( u1_u8_u4_n107 ) , .B2( u1_u8_u4_n143 ) , .A( u1_u8_u4_n174 ) , .B1( u1_u8_u4_n184 ) );
  AOI21_X1 u1_u8_u4_U15 (.B2( u1_u8_u4_n158 ) , .B1( u1_u8_u4_n159 ) , .ZN( u1_u8_u4_n163 ) , .A( u1_u8_u4_n174 ) );
  AOI21_X1 u1_u8_u4_U16 (.A( u1_u8_u4_n153 ) , .B2( u1_u8_u4_n154 ) , .B1( u1_u8_u4_n155 ) , .ZN( u1_u8_u4_n165 ) );
  AOI21_X1 u1_u8_u4_U17 (.A( u1_u8_u4_n156 ) , .B2( u1_u8_u4_n157 ) , .ZN( u1_u8_u4_n164 ) , .B1( u1_u8_u4_n184 ) );
  INV_X1 u1_u8_u4_U18 (.A( u1_u8_u4_n138 ) , .ZN( u1_u8_u4_n170 ) );
  AND2_X1 u1_u8_u4_U19 (.A2( u1_u8_u4_n120 ) , .ZN( u1_u8_u4_n155 ) , .A1( u1_u8_u4_n160 ) );
  INV_X1 u1_u8_u4_U20 (.A( u1_u8_u4_n156 ) , .ZN( u1_u8_u4_n175 ) );
  NAND2_X1 u1_u8_u4_U21 (.A2( u1_u8_u4_n118 ) , .ZN( u1_u8_u4_n131 ) , .A1( u1_u8_u4_n147 ) );
  NAND2_X1 u1_u8_u4_U22 (.A1( u1_u8_u4_n119 ) , .A2( u1_u8_u4_n120 ) , .ZN( u1_u8_u4_n130 ) );
  NAND2_X1 u1_u8_u4_U23 (.ZN( u1_u8_u4_n117 ) , .A2( u1_u8_u4_n118 ) , .A1( u1_u8_u4_n148 ) );
  NAND2_X1 u1_u8_u4_U24 (.ZN( u1_u8_u4_n129 ) , .A1( u1_u8_u4_n134 ) , .A2( u1_u8_u4_n148 ) );
  AND3_X1 u1_u8_u4_U25 (.A1( u1_u8_u4_n119 ) , .A2( u1_u8_u4_n143 ) , .A3( u1_u8_u4_n154 ) , .ZN( u1_u8_u4_n161 ) );
  AND2_X1 u1_u8_u4_U26 (.A1( u1_u8_u4_n145 ) , .A2( u1_u8_u4_n147 ) , .ZN( u1_u8_u4_n159 ) );
  OR3_X1 u1_u8_u4_U27 (.A3( u1_u8_u4_n114 ) , .A2( u1_u8_u4_n115 ) , .A1( u1_u8_u4_n116 ) , .ZN( u1_u8_u4_n136 ) );
  AOI21_X1 u1_u8_u4_U28 (.A( u1_u8_u4_n113 ) , .ZN( u1_u8_u4_n116 ) , .B2( u1_u8_u4_n173 ) , .B1( u1_u8_u4_n174 ) );
  AOI21_X1 u1_u8_u4_U29 (.ZN( u1_u8_u4_n115 ) , .B2( u1_u8_u4_n145 ) , .B1( u1_u8_u4_n146 ) , .A( u1_u8_u4_n156 ) );
  NOR2_X1 u1_u8_u4_U3 (.ZN( u1_u8_u4_n121 ) , .A1( u1_u8_u4_n181 ) , .A2( u1_u8_u4_n182 ) );
  OAI22_X1 u1_u8_u4_U30 (.ZN( u1_u8_u4_n114 ) , .A2( u1_u8_u4_n121 ) , .B1( u1_u8_u4_n160 ) , .B2( u1_u8_u4_n170 ) , .A1( u1_u8_u4_n171 ) );
  INV_X1 u1_u8_u4_U31 (.A( u1_u8_u4_n158 ) , .ZN( u1_u8_u4_n182 ) );
  INV_X1 u1_u8_u4_U32 (.ZN( u1_u8_u4_n181 ) , .A( u1_u8_u4_n96 ) );
  INV_X1 u1_u8_u4_U33 (.A( u1_u8_u4_n144 ) , .ZN( u1_u8_u4_n179 ) );
  INV_X1 u1_u8_u4_U34 (.A( u1_u8_u4_n157 ) , .ZN( u1_u8_u4_n178 ) );
  NAND2_X1 u1_u8_u4_U35 (.A2( u1_u8_u4_n154 ) , .A1( u1_u8_u4_n96 ) , .ZN( u1_u8_u4_n97 ) );
  INV_X1 u1_u8_u4_U36 (.ZN( u1_u8_u4_n186 ) , .A( u1_u8_u4_n95 ) );
  OAI221_X1 u1_u8_u4_U37 (.C1( u1_u8_u4_n134 ) , .B1( u1_u8_u4_n158 ) , .B2( u1_u8_u4_n171 ) , .C2( u1_u8_u4_n173 ) , .A( u1_u8_u4_n94 ) , .ZN( u1_u8_u4_n95 ) );
  AOI222_X1 u1_u8_u4_U38 (.B2( u1_u8_u4_n132 ) , .A1( u1_u8_u4_n138 ) , .C2( u1_u8_u4_n175 ) , .A2( u1_u8_u4_n179 ) , .C1( u1_u8_u4_n181 ) , .B1( u1_u8_u4_n185 ) , .ZN( u1_u8_u4_n94 ) );
  INV_X1 u1_u8_u4_U39 (.A( u1_u8_u4_n113 ) , .ZN( u1_u8_u4_n185 ) );
  INV_X1 u1_u8_u4_U4 (.A( u1_u8_u4_n117 ) , .ZN( u1_u8_u4_n184 ) );
  INV_X1 u1_u8_u4_U40 (.A( u1_u8_u4_n143 ) , .ZN( u1_u8_u4_n183 ) );
  NOR2_X1 u1_u8_u4_U41 (.ZN( u1_u8_u4_n138 ) , .A1( u1_u8_u4_n168 ) , .A2( u1_u8_u4_n169 ) );
  NOR2_X1 u1_u8_u4_U42 (.A1( u1_u8_u4_n150 ) , .A2( u1_u8_u4_n152 ) , .ZN( u1_u8_u4_n153 ) );
  NOR2_X1 u1_u8_u4_U43 (.A2( u1_u8_u4_n128 ) , .A1( u1_u8_u4_n138 ) , .ZN( u1_u8_u4_n156 ) );
  AOI22_X1 u1_u8_u4_U44 (.B2( u1_u8_u4_n122 ) , .A1( u1_u8_u4_n123 ) , .ZN( u1_u8_u4_n124 ) , .B1( u1_u8_u4_n128 ) , .A2( u1_u8_u4_n172 ) );
  INV_X1 u1_u8_u4_U45 (.A( u1_u8_u4_n153 ) , .ZN( u1_u8_u4_n172 ) );
  NAND2_X1 u1_u8_u4_U46 (.A2( u1_u8_u4_n120 ) , .ZN( u1_u8_u4_n123 ) , .A1( u1_u8_u4_n161 ) );
  AOI22_X1 u1_u8_u4_U47 (.B2( u1_u8_u4_n132 ) , .A2( u1_u8_u4_n133 ) , .ZN( u1_u8_u4_n140 ) , .A1( u1_u8_u4_n150 ) , .B1( u1_u8_u4_n179 ) );
  NAND2_X1 u1_u8_u4_U48 (.ZN( u1_u8_u4_n133 ) , .A2( u1_u8_u4_n146 ) , .A1( u1_u8_u4_n154 ) );
  NAND2_X1 u1_u8_u4_U49 (.A1( u1_u8_u4_n103 ) , .ZN( u1_u8_u4_n154 ) , .A2( u1_u8_u4_n98 ) );
  NOR4_X1 u1_u8_u4_U5 (.A4( u1_u8_u4_n106 ) , .A3( u1_u8_u4_n107 ) , .A2( u1_u8_u4_n108 ) , .A1( u1_u8_u4_n109 ) , .ZN( u1_u8_u4_n110 ) );
  NAND2_X1 u1_u8_u4_U50 (.A1( u1_u8_u4_n101 ) , .ZN( u1_u8_u4_n158 ) , .A2( u1_u8_u4_n99 ) );
  AOI21_X1 u1_u8_u4_U51 (.ZN( u1_u8_u4_n127 ) , .A( u1_u8_u4_n136 ) , .B2( u1_u8_u4_n150 ) , .B1( u1_u8_u4_n180 ) );
  INV_X1 u1_u8_u4_U52 (.A( u1_u8_u4_n160 ) , .ZN( u1_u8_u4_n180 ) );
  NAND2_X1 u1_u8_u4_U53 (.A2( u1_u8_u4_n104 ) , .A1( u1_u8_u4_n105 ) , .ZN( u1_u8_u4_n146 ) );
  NAND2_X1 u1_u8_u4_U54 (.A2( u1_u8_u4_n101 ) , .A1( u1_u8_u4_n102 ) , .ZN( u1_u8_u4_n160 ) );
  NAND2_X1 u1_u8_u4_U55 (.ZN( u1_u8_u4_n134 ) , .A1( u1_u8_u4_n98 ) , .A2( u1_u8_u4_n99 ) );
  NAND2_X1 u1_u8_u4_U56 (.A1( u1_u8_u4_n103 ) , .A2( u1_u8_u4_n104 ) , .ZN( u1_u8_u4_n143 ) );
  NAND2_X1 u1_u8_u4_U57 (.A2( u1_u8_u4_n105 ) , .ZN( u1_u8_u4_n145 ) , .A1( u1_u8_u4_n98 ) );
  NAND2_X1 u1_u8_u4_U58 (.A1( u1_u8_u4_n100 ) , .A2( u1_u8_u4_n105 ) , .ZN( u1_u8_u4_n120 ) );
  NAND2_X1 u1_u8_u4_U59 (.A1( u1_u8_u4_n102 ) , .A2( u1_u8_u4_n104 ) , .ZN( u1_u8_u4_n148 ) );
  AOI21_X1 u1_u8_u4_U6 (.ZN( u1_u8_u4_n106 ) , .B2( u1_u8_u4_n146 ) , .B1( u1_u8_u4_n158 ) , .A( u1_u8_u4_n170 ) );
  NAND2_X1 u1_u8_u4_U60 (.A2( u1_u8_u4_n100 ) , .A1( u1_u8_u4_n103 ) , .ZN( u1_u8_u4_n157 ) );
  INV_X1 u1_u8_u4_U61 (.A( u1_u8_u4_n150 ) , .ZN( u1_u8_u4_n173 ) );
  INV_X1 u1_u8_u4_U62 (.A( u1_u8_u4_n152 ) , .ZN( u1_u8_u4_n171 ) );
  NAND2_X1 u1_u8_u4_U63 (.A1( u1_u8_u4_n100 ) , .ZN( u1_u8_u4_n118 ) , .A2( u1_u8_u4_n99 ) );
  NAND2_X1 u1_u8_u4_U64 (.A2( u1_u8_u4_n100 ) , .A1( u1_u8_u4_n102 ) , .ZN( u1_u8_u4_n144 ) );
  NAND2_X1 u1_u8_u4_U65 (.A2( u1_u8_u4_n101 ) , .A1( u1_u8_u4_n105 ) , .ZN( u1_u8_u4_n96 ) );
  INV_X1 u1_u8_u4_U66 (.A( u1_u8_u4_n128 ) , .ZN( u1_u8_u4_n174 ) );
  NAND2_X1 u1_u8_u4_U67 (.A2( u1_u8_u4_n102 ) , .ZN( u1_u8_u4_n119 ) , .A1( u1_u8_u4_n98 ) );
  NAND2_X1 u1_u8_u4_U68 (.A2( u1_u8_u4_n101 ) , .A1( u1_u8_u4_n103 ) , .ZN( u1_u8_u4_n147 ) );
  NAND2_X1 u1_u8_u4_U69 (.A2( u1_u8_u4_n104 ) , .ZN( u1_u8_u4_n113 ) , .A1( u1_u8_u4_n99 ) );
  AOI21_X1 u1_u8_u4_U7 (.ZN( u1_u8_u4_n108 ) , .B2( u1_u8_u4_n134 ) , .B1( u1_u8_u4_n155 ) , .A( u1_u8_u4_n156 ) );
  NOR2_X1 u1_u8_u4_U70 (.A2( u1_u8_X_28 ) , .ZN( u1_u8_u4_n150 ) , .A1( u1_u8_u4_n168 ) );
  NOR2_X1 u1_u8_u4_U71 (.A2( u1_u8_X_29 ) , .ZN( u1_u8_u4_n152 ) , .A1( u1_u8_u4_n169 ) );
  NOR2_X1 u1_u8_u4_U72 (.A2( u1_u8_X_30 ) , .ZN( u1_u8_u4_n105 ) , .A1( u1_u8_u4_n176 ) );
  NOR2_X1 u1_u8_u4_U73 (.A2( u1_u8_X_26 ) , .ZN( u1_u8_u4_n100 ) , .A1( u1_u8_u4_n177 ) );
  NOR2_X1 u1_u8_u4_U74 (.A2( u1_u8_X_28 ) , .A1( u1_u8_X_29 ) , .ZN( u1_u8_u4_n128 ) );
  NOR2_X1 u1_u8_u4_U75 (.A2( u1_u8_X_27 ) , .A1( u1_u8_X_30 ) , .ZN( u1_u8_u4_n102 ) );
  NOR2_X1 u1_u8_u4_U76 (.A2( u1_u8_X_25 ) , .A1( u1_u8_X_26 ) , .ZN( u1_u8_u4_n98 ) );
  AND2_X1 u1_u8_u4_U77 (.A2( u1_u8_X_25 ) , .A1( u1_u8_X_26 ) , .ZN( u1_u8_u4_n104 ) );
  AND2_X1 u1_u8_u4_U78 (.A1( u1_u8_X_30 ) , .A2( u1_u8_u4_n176 ) , .ZN( u1_u8_u4_n99 ) );
  AND2_X1 u1_u8_u4_U79 (.A1( u1_u8_X_26 ) , .ZN( u1_u8_u4_n101 ) , .A2( u1_u8_u4_n177 ) );
  AOI21_X1 u1_u8_u4_U8 (.ZN( u1_u8_u4_n109 ) , .A( u1_u8_u4_n153 ) , .B1( u1_u8_u4_n159 ) , .B2( u1_u8_u4_n184 ) );
  AND2_X1 u1_u8_u4_U80 (.A1( u1_u8_X_27 ) , .A2( u1_u8_X_30 ) , .ZN( u1_u8_u4_n103 ) );
  INV_X1 u1_u8_u4_U81 (.A( u1_u8_X_28 ) , .ZN( u1_u8_u4_n169 ) );
  INV_X1 u1_u8_u4_U82 (.A( u1_u8_X_29 ) , .ZN( u1_u8_u4_n168 ) );
  INV_X1 u1_u8_u4_U83 (.A( u1_u8_X_25 ) , .ZN( u1_u8_u4_n177 ) );
  INV_X1 u1_u8_u4_U84 (.A( u1_u8_X_27 ) , .ZN( u1_u8_u4_n176 ) );
  NAND4_X1 u1_u8_u4_U85 (.ZN( u1_out8_25 ) , .A4( u1_u8_u4_n139 ) , .A3( u1_u8_u4_n140 ) , .A2( u1_u8_u4_n141 ) , .A1( u1_u8_u4_n142 ) );
  OAI21_X1 u1_u8_u4_U86 (.B2( u1_u8_u4_n131 ) , .ZN( u1_u8_u4_n141 ) , .A( u1_u8_u4_n175 ) , .B1( u1_u8_u4_n183 ) );
  OAI21_X1 u1_u8_u4_U87 (.A( u1_u8_u4_n128 ) , .B2( u1_u8_u4_n129 ) , .B1( u1_u8_u4_n130 ) , .ZN( u1_u8_u4_n142 ) );
  NAND4_X1 u1_u8_u4_U88 (.ZN( u1_out8_14 ) , .A4( u1_u8_u4_n124 ) , .A3( u1_u8_u4_n125 ) , .A2( u1_u8_u4_n126 ) , .A1( u1_u8_u4_n127 ) );
  AOI22_X1 u1_u8_u4_U89 (.B2( u1_u8_u4_n117 ) , .ZN( u1_u8_u4_n126 ) , .A1( u1_u8_u4_n129 ) , .B1( u1_u8_u4_n152 ) , .A2( u1_u8_u4_n175 ) );
  AOI211_X1 u1_u8_u4_U9 (.B( u1_u8_u4_n136 ) , .A( u1_u8_u4_n137 ) , .C2( u1_u8_u4_n138 ) , .ZN( u1_u8_u4_n139 ) , .C1( u1_u8_u4_n182 ) );
  AOI22_X1 u1_u8_u4_U90 (.ZN( u1_u8_u4_n125 ) , .B2( u1_u8_u4_n131 ) , .A2( u1_u8_u4_n132 ) , .B1( u1_u8_u4_n138 ) , .A1( u1_u8_u4_n178 ) );
  NAND4_X1 u1_u8_u4_U91 (.ZN( u1_out8_8 ) , .A4( u1_u8_u4_n110 ) , .A3( u1_u8_u4_n111 ) , .A2( u1_u8_u4_n112 ) , .A1( u1_u8_u4_n186 ) );
  NAND2_X1 u1_u8_u4_U92 (.ZN( u1_u8_u4_n112 ) , .A2( u1_u8_u4_n130 ) , .A1( u1_u8_u4_n150 ) );
  AOI22_X1 u1_u8_u4_U93 (.ZN( u1_u8_u4_n111 ) , .B2( u1_u8_u4_n132 ) , .A1( u1_u8_u4_n152 ) , .B1( u1_u8_u4_n178 ) , .A2( u1_u8_u4_n97 ) );
  AOI22_X1 u1_u8_u4_U94 (.B2( u1_u8_u4_n149 ) , .B1( u1_u8_u4_n150 ) , .A2( u1_u8_u4_n151 ) , .A1( u1_u8_u4_n152 ) , .ZN( u1_u8_u4_n167 ) );
  NOR4_X1 u1_u8_u4_U95 (.A4( u1_u8_u4_n162 ) , .A3( u1_u8_u4_n163 ) , .A2( u1_u8_u4_n164 ) , .A1( u1_u8_u4_n165 ) , .ZN( u1_u8_u4_n166 ) );
  NAND3_X1 u1_u8_u4_U96 (.ZN( u1_out8_3 ) , .A3( u1_u8_u4_n166 ) , .A1( u1_u8_u4_n167 ) , .A2( u1_u8_u4_n186 ) );
  NAND3_X1 u1_u8_u4_U97 (.A3( u1_u8_u4_n146 ) , .A2( u1_u8_u4_n147 ) , .A1( u1_u8_u4_n148 ) , .ZN( u1_u8_u4_n149 ) );
  NAND3_X1 u1_u8_u4_U98 (.A3( u1_u8_u4_n143 ) , .A2( u1_u8_u4_n144 ) , .A1( u1_u8_u4_n145 ) , .ZN( u1_u8_u4_n151 ) );
  NAND3_X1 u1_u8_u4_U99 (.A3( u1_u8_u4_n121 ) , .ZN( u1_u8_u4_n122 ) , .A2( u1_u8_u4_n144 ) , .A1( u1_u8_u4_n154 ) );
  XOR2_X1 u1_u9_U26 (.B( u1_K10_30 ) , .A( u1_R8_21 ) , .Z( u1_u9_X_30 ) );
  XOR2_X1 u1_u9_U28 (.B( u1_K10_29 ) , .A( u1_R8_20 ) , .Z( u1_u9_X_29 ) );
  XOR2_X1 u1_u9_U29 (.B( u1_K10_28 ) , .A( u1_R8_19 ) , .Z( u1_u9_X_28 ) );
  XOR2_X1 u1_u9_U30 (.B( u1_K10_27 ) , .A( u1_R8_18 ) , .Z( u1_u9_X_27 ) );
  XOR2_X1 u1_u9_U31 (.B( u1_K10_26 ) , .A( u1_R8_17 ) , .Z( u1_u9_X_26 ) );
  XOR2_X1 u1_u9_U32 (.B( u1_K10_25 ) , .A( u1_R8_16 ) , .Z( u1_u9_X_25 ) );
  OAI22_X1 u1_u9_u4_U10 (.B2( u1_u9_u4_n135 ) , .ZN( u1_u9_u4_n137 ) , .B1( u1_u9_u4_n153 ) , .A1( u1_u9_u4_n155 ) , .A2( u1_u9_u4_n171 ) );
  AND3_X1 u1_u9_u4_U11 (.A2( u1_u9_u4_n134 ) , .ZN( u1_u9_u4_n135 ) , .A3( u1_u9_u4_n145 ) , .A1( u1_u9_u4_n157 ) );
  NAND2_X1 u1_u9_u4_U12 (.ZN( u1_u9_u4_n132 ) , .A2( u1_u9_u4_n170 ) , .A1( u1_u9_u4_n173 ) );
  AOI21_X1 u1_u9_u4_U13 (.B2( u1_u9_u4_n160 ) , .B1( u1_u9_u4_n161 ) , .ZN( u1_u9_u4_n162 ) , .A( u1_u9_u4_n170 ) );
  AOI21_X1 u1_u9_u4_U14 (.ZN( u1_u9_u4_n107 ) , .B2( u1_u9_u4_n143 ) , .A( u1_u9_u4_n174 ) , .B1( u1_u9_u4_n184 ) );
  AOI21_X1 u1_u9_u4_U15 (.B2( u1_u9_u4_n158 ) , .B1( u1_u9_u4_n159 ) , .ZN( u1_u9_u4_n163 ) , .A( u1_u9_u4_n174 ) );
  AOI21_X1 u1_u9_u4_U16 (.A( u1_u9_u4_n153 ) , .B2( u1_u9_u4_n154 ) , .B1( u1_u9_u4_n155 ) , .ZN( u1_u9_u4_n165 ) );
  AOI21_X1 u1_u9_u4_U17 (.A( u1_u9_u4_n156 ) , .B2( u1_u9_u4_n157 ) , .ZN( u1_u9_u4_n164 ) , .B1( u1_u9_u4_n184 ) );
  INV_X1 u1_u9_u4_U18 (.A( u1_u9_u4_n138 ) , .ZN( u1_u9_u4_n170 ) );
  AND2_X1 u1_u9_u4_U19 (.A2( u1_u9_u4_n120 ) , .ZN( u1_u9_u4_n155 ) , .A1( u1_u9_u4_n160 ) );
  INV_X1 u1_u9_u4_U20 (.A( u1_u9_u4_n156 ) , .ZN( u1_u9_u4_n175 ) );
  NAND2_X1 u1_u9_u4_U21 (.A2( u1_u9_u4_n118 ) , .ZN( u1_u9_u4_n131 ) , .A1( u1_u9_u4_n147 ) );
  NAND2_X1 u1_u9_u4_U22 (.A1( u1_u9_u4_n119 ) , .A2( u1_u9_u4_n120 ) , .ZN( u1_u9_u4_n130 ) );
  NAND2_X1 u1_u9_u4_U23 (.ZN( u1_u9_u4_n117 ) , .A2( u1_u9_u4_n118 ) , .A1( u1_u9_u4_n148 ) );
  NAND2_X1 u1_u9_u4_U24 (.ZN( u1_u9_u4_n129 ) , .A1( u1_u9_u4_n134 ) , .A2( u1_u9_u4_n148 ) );
  AND3_X1 u1_u9_u4_U25 (.A1( u1_u9_u4_n119 ) , .A2( u1_u9_u4_n143 ) , .A3( u1_u9_u4_n154 ) , .ZN( u1_u9_u4_n161 ) );
  AND2_X1 u1_u9_u4_U26 (.A1( u1_u9_u4_n145 ) , .A2( u1_u9_u4_n147 ) , .ZN( u1_u9_u4_n159 ) );
  OR3_X1 u1_u9_u4_U27 (.A3( u1_u9_u4_n114 ) , .A2( u1_u9_u4_n115 ) , .A1( u1_u9_u4_n116 ) , .ZN( u1_u9_u4_n136 ) );
  AOI21_X1 u1_u9_u4_U28 (.A( u1_u9_u4_n113 ) , .ZN( u1_u9_u4_n116 ) , .B2( u1_u9_u4_n173 ) , .B1( u1_u9_u4_n174 ) );
  AOI21_X1 u1_u9_u4_U29 (.ZN( u1_u9_u4_n115 ) , .B2( u1_u9_u4_n145 ) , .B1( u1_u9_u4_n146 ) , .A( u1_u9_u4_n156 ) );
  NOR2_X1 u1_u9_u4_U3 (.ZN( u1_u9_u4_n121 ) , .A1( u1_u9_u4_n181 ) , .A2( u1_u9_u4_n182 ) );
  OAI22_X1 u1_u9_u4_U30 (.ZN( u1_u9_u4_n114 ) , .A2( u1_u9_u4_n121 ) , .B1( u1_u9_u4_n160 ) , .B2( u1_u9_u4_n170 ) , .A1( u1_u9_u4_n171 ) );
  INV_X1 u1_u9_u4_U31 (.A( u1_u9_u4_n158 ) , .ZN( u1_u9_u4_n182 ) );
  INV_X1 u1_u9_u4_U32 (.ZN( u1_u9_u4_n181 ) , .A( u1_u9_u4_n96 ) );
  INV_X1 u1_u9_u4_U33 (.A( u1_u9_u4_n144 ) , .ZN( u1_u9_u4_n179 ) );
  INV_X1 u1_u9_u4_U34 (.A( u1_u9_u4_n157 ) , .ZN( u1_u9_u4_n178 ) );
  NAND2_X1 u1_u9_u4_U35 (.A2( u1_u9_u4_n154 ) , .A1( u1_u9_u4_n96 ) , .ZN( u1_u9_u4_n97 ) );
  INV_X1 u1_u9_u4_U36 (.ZN( u1_u9_u4_n186 ) , .A( u1_u9_u4_n95 ) );
  OAI221_X1 u1_u9_u4_U37 (.C1( u1_u9_u4_n134 ) , .B1( u1_u9_u4_n158 ) , .B2( u1_u9_u4_n171 ) , .C2( u1_u9_u4_n173 ) , .A( u1_u9_u4_n94 ) , .ZN( u1_u9_u4_n95 ) );
  AOI222_X1 u1_u9_u4_U38 (.B2( u1_u9_u4_n132 ) , .A1( u1_u9_u4_n138 ) , .C2( u1_u9_u4_n175 ) , .A2( u1_u9_u4_n179 ) , .C1( u1_u9_u4_n181 ) , .B1( u1_u9_u4_n185 ) , .ZN( u1_u9_u4_n94 ) );
  INV_X1 u1_u9_u4_U39 (.A( u1_u9_u4_n113 ) , .ZN( u1_u9_u4_n185 ) );
  INV_X1 u1_u9_u4_U4 (.A( u1_u9_u4_n117 ) , .ZN( u1_u9_u4_n184 ) );
  INV_X1 u1_u9_u4_U40 (.A( u1_u9_u4_n143 ) , .ZN( u1_u9_u4_n183 ) );
  NOR2_X1 u1_u9_u4_U41 (.ZN( u1_u9_u4_n138 ) , .A1( u1_u9_u4_n168 ) , .A2( u1_u9_u4_n169 ) );
  NOR2_X1 u1_u9_u4_U42 (.A1( u1_u9_u4_n150 ) , .A2( u1_u9_u4_n152 ) , .ZN( u1_u9_u4_n153 ) );
  NOR2_X1 u1_u9_u4_U43 (.A2( u1_u9_u4_n128 ) , .A1( u1_u9_u4_n138 ) , .ZN( u1_u9_u4_n156 ) );
  AOI22_X1 u1_u9_u4_U44 (.B2( u1_u9_u4_n122 ) , .A1( u1_u9_u4_n123 ) , .ZN( u1_u9_u4_n124 ) , .B1( u1_u9_u4_n128 ) , .A2( u1_u9_u4_n172 ) );
  INV_X1 u1_u9_u4_U45 (.A( u1_u9_u4_n153 ) , .ZN( u1_u9_u4_n172 ) );
  NAND2_X1 u1_u9_u4_U46 (.A2( u1_u9_u4_n120 ) , .ZN( u1_u9_u4_n123 ) , .A1( u1_u9_u4_n161 ) );
  AOI22_X1 u1_u9_u4_U47 (.B2( u1_u9_u4_n132 ) , .A2( u1_u9_u4_n133 ) , .ZN( u1_u9_u4_n140 ) , .A1( u1_u9_u4_n150 ) , .B1( u1_u9_u4_n179 ) );
  NAND2_X1 u1_u9_u4_U48 (.ZN( u1_u9_u4_n133 ) , .A2( u1_u9_u4_n146 ) , .A1( u1_u9_u4_n154 ) );
  NAND2_X1 u1_u9_u4_U49 (.A1( u1_u9_u4_n103 ) , .ZN( u1_u9_u4_n154 ) , .A2( u1_u9_u4_n98 ) );
  NOR4_X1 u1_u9_u4_U5 (.A4( u1_u9_u4_n106 ) , .A3( u1_u9_u4_n107 ) , .A2( u1_u9_u4_n108 ) , .A1( u1_u9_u4_n109 ) , .ZN( u1_u9_u4_n110 ) );
  NAND2_X1 u1_u9_u4_U50 (.A1( u1_u9_u4_n101 ) , .ZN( u1_u9_u4_n158 ) , .A2( u1_u9_u4_n99 ) );
  AOI21_X1 u1_u9_u4_U51 (.ZN( u1_u9_u4_n127 ) , .A( u1_u9_u4_n136 ) , .B2( u1_u9_u4_n150 ) , .B1( u1_u9_u4_n180 ) );
  INV_X1 u1_u9_u4_U52 (.A( u1_u9_u4_n160 ) , .ZN( u1_u9_u4_n180 ) );
  NAND2_X1 u1_u9_u4_U53 (.A2( u1_u9_u4_n104 ) , .A1( u1_u9_u4_n105 ) , .ZN( u1_u9_u4_n146 ) );
  NAND2_X1 u1_u9_u4_U54 (.A2( u1_u9_u4_n101 ) , .A1( u1_u9_u4_n102 ) , .ZN( u1_u9_u4_n160 ) );
  NAND2_X1 u1_u9_u4_U55 (.ZN( u1_u9_u4_n134 ) , .A1( u1_u9_u4_n98 ) , .A2( u1_u9_u4_n99 ) );
  NAND2_X1 u1_u9_u4_U56 (.A1( u1_u9_u4_n103 ) , .A2( u1_u9_u4_n104 ) , .ZN( u1_u9_u4_n143 ) );
  NAND2_X1 u1_u9_u4_U57 (.A2( u1_u9_u4_n105 ) , .ZN( u1_u9_u4_n145 ) , .A1( u1_u9_u4_n98 ) );
  NAND2_X1 u1_u9_u4_U58 (.A1( u1_u9_u4_n100 ) , .A2( u1_u9_u4_n105 ) , .ZN( u1_u9_u4_n120 ) );
  NAND2_X1 u1_u9_u4_U59 (.A1( u1_u9_u4_n102 ) , .A2( u1_u9_u4_n104 ) , .ZN( u1_u9_u4_n148 ) );
  AOI21_X1 u1_u9_u4_U6 (.ZN( u1_u9_u4_n106 ) , .B2( u1_u9_u4_n146 ) , .B1( u1_u9_u4_n158 ) , .A( u1_u9_u4_n170 ) );
  NAND2_X1 u1_u9_u4_U60 (.A2( u1_u9_u4_n100 ) , .A1( u1_u9_u4_n103 ) , .ZN( u1_u9_u4_n157 ) );
  INV_X1 u1_u9_u4_U61 (.A( u1_u9_u4_n150 ) , .ZN( u1_u9_u4_n173 ) );
  INV_X1 u1_u9_u4_U62 (.A( u1_u9_u4_n152 ) , .ZN( u1_u9_u4_n171 ) );
  NAND2_X1 u1_u9_u4_U63 (.A1( u1_u9_u4_n100 ) , .ZN( u1_u9_u4_n118 ) , .A2( u1_u9_u4_n99 ) );
  NAND2_X1 u1_u9_u4_U64 (.A2( u1_u9_u4_n100 ) , .A1( u1_u9_u4_n102 ) , .ZN( u1_u9_u4_n144 ) );
  NAND2_X1 u1_u9_u4_U65 (.A2( u1_u9_u4_n101 ) , .A1( u1_u9_u4_n105 ) , .ZN( u1_u9_u4_n96 ) );
  INV_X1 u1_u9_u4_U66 (.A( u1_u9_u4_n128 ) , .ZN( u1_u9_u4_n174 ) );
  NAND2_X1 u1_u9_u4_U67 (.A2( u1_u9_u4_n102 ) , .ZN( u1_u9_u4_n119 ) , .A1( u1_u9_u4_n98 ) );
  NAND2_X1 u1_u9_u4_U68 (.A2( u1_u9_u4_n101 ) , .A1( u1_u9_u4_n103 ) , .ZN( u1_u9_u4_n147 ) );
  NAND2_X1 u1_u9_u4_U69 (.A2( u1_u9_u4_n104 ) , .ZN( u1_u9_u4_n113 ) , .A1( u1_u9_u4_n99 ) );
  AOI21_X1 u1_u9_u4_U7 (.ZN( u1_u9_u4_n108 ) , .B2( u1_u9_u4_n134 ) , .B1( u1_u9_u4_n155 ) , .A( u1_u9_u4_n156 ) );
  NOR2_X1 u1_u9_u4_U70 (.A2( u1_u9_X_28 ) , .ZN( u1_u9_u4_n150 ) , .A1( u1_u9_u4_n168 ) );
  NOR2_X1 u1_u9_u4_U71 (.A2( u1_u9_X_29 ) , .ZN( u1_u9_u4_n152 ) , .A1( u1_u9_u4_n169 ) );
  NOR2_X1 u1_u9_u4_U72 (.A2( u1_u9_X_30 ) , .ZN( u1_u9_u4_n105 ) , .A1( u1_u9_u4_n176 ) );
  NOR2_X1 u1_u9_u4_U73 (.A2( u1_u9_X_26 ) , .ZN( u1_u9_u4_n100 ) , .A1( u1_u9_u4_n177 ) );
  NOR2_X1 u1_u9_u4_U74 (.A2( u1_u9_X_28 ) , .A1( u1_u9_X_29 ) , .ZN( u1_u9_u4_n128 ) );
  NOR2_X1 u1_u9_u4_U75 (.A2( u1_u9_X_27 ) , .A1( u1_u9_X_30 ) , .ZN( u1_u9_u4_n102 ) );
  NOR2_X1 u1_u9_u4_U76 (.A2( u1_u9_X_25 ) , .A1( u1_u9_X_26 ) , .ZN( u1_u9_u4_n98 ) );
  AND2_X1 u1_u9_u4_U77 (.A2( u1_u9_X_25 ) , .A1( u1_u9_X_26 ) , .ZN( u1_u9_u4_n104 ) );
  AND2_X1 u1_u9_u4_U78 (.A1( u1_u9_X_30 ) , .A2( u1_u9_u4_n176 ) , .ZN( u1_u9_u4_n99 ) );
  AND2_X1 u1_u9_u4_U79 (.A1( u1_u9_X_26 ) , .ZN( u1_u9_u4_n101 ) , .A2( u1_u9_u4_n177 ) );
  AOI21_X1 u1_u9_u4_U8 (.ZN( u1_u9_u4_n109 ) , .A( u1_u9_u4_n153 ) , .B1( u1_u9_u4_n159 ) , .B2( u1_u9_u4_n184 ) );
  AND2_X1 u1_u9_u4_U80 (.A1( u1_u9_X_27 ) , .A2( u1_u9_X_30 ) , .ZN( u1_u9_u4_n103 ) );
  INV_X1 u1_u9_u4_U81 (.A( u1_u9_X_28 ) , .ZN( u1_u9_u4_n169 ) );
  INV_X1 u1_u9_u4_U82 (.A( u1_u9_X_29 ) , .ZN( u1_u9_u4_n168 ) );
  INV_X1 u1_u9_u4_U83 (.A( u1_u9_X_25 ) , .ZN( u1_u9_u4_n177 ) );
  INV_X1 u1_u9_u4_U84 (.A( u1_u9_X_27 ) , .ZN( u1_u9_u4_n176 ) );
  NAND4_X1 u1_u9_u4_U85 (.ZN( u1_out9_25 ) , .A4( u1_u9_u4_n139 ) , .A3( u1_u9_u4_n140 ) , .A2( u1_u9_u4_n141 ) , .A1( u1_u9_u4_n142 ) );
  OAI21_X1 u1_u9_u4_U86 (.A( u1_u9_u4_n128 ) , .B2( u1_u9_u4_n129 ) , .B1( u1_u9_u4_n130 ) , .ZN( u1_u9_u4_n142 ) );
  OAI21_X1 u1_u9_u4_U87 (.B2( u1_u9_u4_n131 ) , .ZN( u1_u9_u4_n141 ) , .A( u1_u9_u4_n175 ) , .B1( u1_u9_u4_n183 ) );
  NAND4_X1 u1_u9_u4_U88 (.ZN( u1_out9_14 ) , .A4( u1_u9_u4_n124 ) , .A3( u1_u9_u4_n125 ) , .A2( u1_u9_u4_n126 ) , .A1( u1_u9_u4_n127 ) );
  AOI22_X1 u1_u9_u4_U89 (.B2( u1_u9_u4_n117 ) , .ZN( u1_u9_u4_n126 ) , .A1( u1_u9_u4_n129 ) , .B1( u1_u9_u4_n152 ) , .A2( u1_u9_u4_n175 ) );
  AOI211_X1 u1_u9_u4_U9 (.B( u1_u9_u4_n136 ) , .A( u1_u9_u4_n137 ) , .C2( u1_u9_u4_n138 ) , .ZN( u1_u9_u4_n139 ) , .C1( u1_u9_u4_n182 ) );
  AOI22_X1 u1_u9_u4_U90 (.ZN( u1_u9_u4_n125 ) , .B2( u1_u9_u4_n131 ) , .A2( u1_u9_u4_n132 ) , .B1( u1_u9_u4_n138 ) , .A1( u1_u9_u4_n178 ) );
  NAND4_X1 u1_u9_u4_U91 (.ZN( u1_out9_8 ) , .A4( u1_u9_u4_n110 ) , .A3( u1_u9_u4_n111 ) , .A2( u1_u9_u4_n112 ) , .A1( u1_u9_u4_n186 ) );
  NAND2_X1 u1_u9_u4_U92 (.ZN( u1_u9_u4_n112 ) , .A2( u1_u9_u4_n130 ) , .A1( u1_u9_u4_n150 ) );
  AOI22_X1 u1_u9_u4_U93 (.ZN( u1_u9_u4_n111 ) , .B2( u1_u9_u4_n132 ) , .A1( u1_u9_u4_n152 ) , .B1( u1_u9_u4_n178 ) , .A2( u1_u9_u4_n97 ) );
  AOI22_X1 u1_u9_u4_U94 (.B2( u1_u9_u4_n149 ) , .B1( u1_u9_u4_n150 ) , .A2( u1_u9_u4_n151 ) , .A1( u1_u9_u4_n152 ) , .ZN( u1_u9_u4_n167 ) );
  NOR4_X1 u1_u9_u4_U95 (.A4( u1_u9_u4_n162 ) , .A3( u1_u9_u4_n163 ) , .A2( u1_u9_u4_n164 ) , .A1( u1_u9_u4_n165 ) , .ZN( u1_u9_u4_n166 ) );
  NAND3_X1 u1_u9_u4_U96 (.ZN( u1_out9_3 ) , .A3( u1_u9_u4_n166 ) , .A1( u1_u9_u4_n167 ) , .A2( u1_u9_u4_n186 ) );
  NAND3_X1 u1_u9_u4_U97 (.A3( u1_u9_u4_n146 ) , .A2( u1_u9_u4_n147 ) , .A1( u1_u9_u4_n148 ) , .ZN( u1_u9_u4_n149 ) );
  NAND3_X1 u1_u9_u4_U98 (.A3( u1_u9_u4_n143 ) , .A2( u1_u9_u4_n144 ) , .A1( u1_u9_u4_n145 ) , .ZN( u1_u9_u4_n151 ) );
  NAND3_X1 u1_u9_u4_U99 (.A3( u1_u9_u4_n121 ) , .ZN( u1_u9_u4_n122 ) , .A2( u1_u9_u4_n144 ) , .A1( u1_u9_u4_n154 ) );
  AOI22_X1 u1_uk_U100 (.B2( u1_uk_K_r0_28 ) , .A2( u1_uk_K_r0_49 ) , .ZN( u1_uk_n1031 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U1010 (.ZN( u1_K5_4 ) , .A( u1_uk_n1085 ) , .B2( u1_uk_n1411 ) , .B1( u1_uk_n60 ) );
  NAND2_X1 u1_uk_U1011 (.A1( u1_uk_K_r3_4 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1085 ) );
  OAI21_X1 u1_uk_U1014 (.ZN( u1_K3_5 ) , .B1( u1_uk_n102 ) , .A( u1_uk_n1048 ) , .B2( u1_uk_n1332 ) );
  NAND2_X1 u1_uk_U1015 (.A1( u1_uk_K_r1_10 ) , .ZN( u1_uk_n1048 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U102 (.ZN( u1_K13_41 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1753 ) , .A2( u1_uk_n1768 ) , .A1( u1_uk_n209 ) );
  OAI21_X1 u1_uk_U1050 (.ZN( u1_K8_28 ) , .A( u1_uk_n1133 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1562 ) );
  NAND2_X1 u1_uk_U1051 (.A1( u1_uk_K_r6_51 ) , .ZN( u1_uk_n1133 ) , .A2( u1_uk_n145 ) );
  OAI21_X1 u1_uk_U1056 (.ZN( u1_K7_31 ) , .A( u1_uk_n1117 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1508 ) );
  NAND2_X1 u1_uk_U1057 (.A1( u1_uk_K_r5_16 ) , .ZN( u1_uk_n1117 ) , .A2( u1_uk_n17 ) );
  INV_X1 u1_uk_U1153 (.ZN( u1_K7_32 ) , .A( u1_uk_n1118 ) );
  AOI22_X1 u1_uk_U1154 (.B2( u1_uk_K_r5_0 ) , .A2( u1_uk_K_r5_51 ) , .ZN( u1_uk_n1118 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n222 ) );
  OAI22_X1 u1_uk_U116 (.ZN( u1_K7_5 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1487 ) , .A2( u1_uk_n1504 ) , .B1( u1_uk_n242 ) );
  OAI22_X1 u1_uk_U117 (.ZN( u1_K5_5 ) , .A1( u1_uk_n128 ) , .A2( u1_uk_n1398 ) , .B2( u1_uk_n1422 ) , .B1( u1_uk_n242 ) );
  INV_X1 u1_uk_U12 (.A( u1_uk_n208 ) , .ZN( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U124 (.ZN( u1_K13_47 ) , .A1( u1_uk_n117 ) , .B2( u1_uk_n1782 ) , .A2( u1_uk_n1792 ) , .B1( u1_uk_n208 ) );
  INV_X1 u1_uk_U13 (.A( u1_uk_n222 ) , .ZN( u1_uk_n99 ) );
  OAI21_X1 u1_uk_U139 (.ZN( u1_K5_15 ) , .A( u1_uk_n1072 ) , .B2( u1_uk_n1409 ) , .B1( u1_uk_n93 ) );
  NAND2_X1 u1_uk_U140 (.A1( u1_uk_K_r3_34 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1072 ) );
  INV_X1 u1_uk_U141 (.ZN( u1_K13_15 ) , .A( u1_uk_n678 ) );
  AOI22_X1 u1_uk_U142 (.B2( u1_uk_K_r11_11 ) , .A2( u1_uk_K_r11_48 ) , .B1( u1_uk_n162 ) , .A1( u1_uk_n240 ) , .ZN( u1_uk_n678 ) );
  OAI22_X1 u1_uk_U146 (.ZN( u1_K3_15 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1312 ) , .B2( u1_uk_n1347 ) , .A1( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U167 (.ZN( u1_K3_19 ) , .A( u1_uk_n1037 ) , .B2( u1_uk_n1324 ) , .B1( u1_uk_n155 ) );
  NAND2_X1 u1_uk_U168 (.A1( u1_uk_K_r1_33 ) , .ZN( u1_uk_n1037 ) , .A2( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U175 (.ZN( u1_K2_30 ) , .B2( u1_uk_n1260 ) , .A2( u1_uk_n1289 ) , .A1( u1_uk_n257 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U176 (.ZN( u1_K14_30 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1811 ) , .A2( u1_uk_n1838 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U179 (.ZN( u1_K10_30 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1628 ) , .A2( u1_uk_n1656 ) , .B1( u1_uk_n250 ) );
  OAI21_X1 u1_uk_U184 (.ZN( u1_K8_30 ) , .A( u1_uk_n1136 ) , .B2( u1_uk_n1555 ) , .B1( u1_uk_n207 ) );
  NAND2_X1 u1_uk_U185 (.A1( u1_uk_K_r6_29 ) , .ZN( u1_uk_n1136 ) , .A2( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U188 (.ZN( u1_K13_14 ) , .A1( u1_uk_n147 ) , .B2( u1_uk_n1756 ) , .A2( u1_uk_n1780 ) , .B1( u1_uk_n203 ) );
  INV_X1 u1_uk_U19 (.ZN( u1_uk_n141 ) , .A( u1_uk_n238 ) );
  INV_X1 u1_uk_U206 (.ZN( u1_K3_24 ) , .A( u1_uk_n1038 ) );
  AOI22_X1 u1_uk_U207 (.B2( u1_uk_K_r1_17 ) , .A2( u1_uk_K_r1_41 ) , .ZN( u1_uk_n1038 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n294 ) );
  OAI21_X1 u1_uk_U211 (.ZN( u1_K9_30 ) , .A( u1_uk_n1161 ) , .B2( u1_uk_n1600 ) , .B1( u1_uk_n27 ) );
  NAND2_X1 u1_uk_U212 (.A1( u1_uk_K_r7_29 ) , .ZN( u1_uk_n1161 ) , .A2( u1_uk_n187 ) );
  OAI22_X1 u1_uk_U217 (.ZN( u1_K3_14 ) , .B2( u1_uk_n1340 ) , .A2( u1_uk_n1347 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n31 ) );
  INV_X1 u1_uk_U22 (.ZN( u1_uk_n147 ) , .A( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U223 (.ZN( u1_K8_31 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1529 ) , .A2( u1_uk_n1567 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U244 (.ZN( u1_K14_31 ) , .A1( u1_uk_n109 ) , .B2( u1_uk_n1827 ) , .A2( u1_uk_n1833 ) , .B1( u1_uk_n223 ) );
  OAI22_X1 u1_uk_U248 (.ZN( u1_K13_39 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1755 ) , .A2( u1_uk_n1774 ) , .B1( u1_uk_n240 ) );
  INV_X1 u1_uk_U26 (.ZN( u1_uk_n145 ) , .A( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U267 (.ZN( u1_K13_44 ) , .B2( u1_uk_n1754 ) , .A2( u1_uk_n1769 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n31 ) );
  OAI21_X1 u1_uk_U268 (.ZN( u1_K13_48 ) , .B1( u1_uk_n129 ) , .B2( u1_uk_n1785 ) , .A( u1_uk_n947 ) );
  NAND2_X1 u1_uk_U269 (.A1( u1_uk_K_r11_8 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n947 ) );
  INV_X1 u1_uk_U27 (.ZN( u1_uk_n148 ) , .A( u1_uk_n214 ) );
  INV_X1 u1_uk_U28 (.A( u1_uk_n202 ) , .ZN( u1_uk_n27 ) );
  INV_X1 u1_uk_U29 (.ZN( u1_uk_n10 ) , .A( u1_uk_n220 ) );
  OAI21_X1 u1_uk_U293 (.ZN( u1_K5_6 ) , .A( u1_uk_n1086 ) , .B2( u1_uk_n1417 ) , .B1( u1_uk_n93 ) );
  NAND2_X1 u1_uk_U294 (.A1( u1_uk_K_r3_10 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n1086 ) );
  INV_X1 u1_uk_U3 (.A( u1_uk_n191 ) , .ZN( u1_uk_n31 ) );
  INV_X1 u1_uk_U30 (.ZN( u1_uk_n17 ) , .A( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U308 (.ZN( u1_K3_8 ) , .A2( u1_uk_n1310 ) , .B2( u1_uk_n1326 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n94 ) );
  INV_X1 u1_uk_U31 (.ZN( u1_uk_n11 ) , .A( u1_uk_n217 ) );
  INV_X1 u1_uk_U315 (.ZN( u1_K9_26 ) , .A( u1_uk_n1158 ) );
  AOI22_X1 u1_uk_U316 (.B2( u1_uk_K_r7_15 ) , .A2( u1_uk_K_r7_8 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1158 ) , .B1( u1_uk_n208 ) );
  INV_X1 u1_uk_U32 (.ZN( u1_uk_n155 ) , .A( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U328 (.ZN( u1_K2_26 ) , .B2( u1_uk_n1289 ) , .A2( u1_uk_n1295 ) , .A1( u1_uk_n214 ) , .B1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U330 (.ZN( u1_K14_26 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1822 ) , .A2( u1_uk_n1839 ) , .A1( u1_uk_n209 ) );
  OAI22_X1 u1_uk_U332 (.ZN( u1_K10_26 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1639 ) , .A2( u1_uk_n1655 ) , .A1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U333 (.ZN( u1_K8_26 ) , .A1( u1_uk_n10 ) , .A2( u1_uk_n1533 ) , .B2( u1_uk_n1540 ) , .B1( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U337 (.ZN( u1_K13_46 ) , .B1( u1_uk_n147 ) , .B2( u1_uk_n1763 ) , .A2( u1_uk_n1775 ) , .A1( u1_uk_n214 ) );
  INV_X1 u1_uk_U34 (.ZN( u1_uk_n162 ) , .A( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U348 (.ZN( u1_K7_4 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1504 ) , .A2( u1_uk_n1527 ) , .B1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U355 (.ZN( u1_K3_4 ) , .B2( u1_uk_n1323 ) , .A2( u1_uk_n1331 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n94 ) );
  OAI22_X1 u1_uk_U363 (.ZN( u1_K13_40 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1774 ) , .A2( u1_uk_n1784 ) , .B1( u1_uk_n252 ) );
  OAI22_X1 u1_uk_U377 (.ZN( u1_K2_40 ) , .A2( u1_uk_n1265 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1296 ) , .B1( u1_uk_n223 ) );
  BUF_X1 u1_uk_U38 (.Z( u1_uk_n208 ) , .A( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U384 (.ZN( u1_K14_28 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1821 ) , .A2( u1_uk_n1827 ) , .B1( u1_uk_n222 ) );
  BUF_X1 u1_uk_U39 (.Z( u1_uk_n202 ) , .A( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U392 (.ZN( u1_K10_28 ) , .A1( u1_uk_n128 ) , .B2( u1_uk_n1640 ) , .A2( u1_uk_n1647 ) , .B1( u1_uk_n240 ) );
  OAI22_X1 u1_uk_U393 (.ZN( u1_K9_28 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1607 ) , .A2( u1_uk_n1614 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U398 (.ZN( u1_K3_1 ) , .B2( u1_uk_n1315 ) , .A2( u1_uk_n1320 ) , .A1( u1_uk_n279 ) , .B1( u1_uk_n83 ) );
  BUF_X1 u1_uk_U40 (.Z( u1_uk_n209 ) , .A( u1_uk_n286 ) );
  OAI21_X1 u1_uk_U400 (.ZN( u1_K7_1 ) , .A( u1_uk_n1108 ) , .B2( u1_uk_n1492 ) , .B1( u1_uk_n217 ) );
  NAND2_X1 u1_uk_U401 (.A1( u1_uk_K_r5_10 ) , .ZN( u1_uk_n1108 ) , .A2( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U402 (.ZN( u1_K5_1 ) , .B2( u1_uk_n1422 ) , .A2( u1_uk_n1429 ) , .B1( u1_uk_n164 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U404 (.ZN( u1_K13_16 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1761 ) , .A2( u1_uk_n1766 ) , .B1( u1_uk_n202 ) );
  OAI21_X1 u1_uk_U413 (.ZN( u1_K3_16 ) , .A( u1_uk_n1036 ) , .B2( u1_uk_n1348 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U414 (.A1( u1_uk_K_r1_6 ) , .ZN( u1_uk_n1036 ) , .A2( u1_uk_n99 ) );
  BUF_X1 u1_uk_U42 (.Z( u1_uk_n242 ) , .A( u1_uk_n271 ) );
  OAI21_X1 u1_uk_U426 (.ZN( u1_K3_9 ) , .A( u1_uk_n1049 ) , .B2( u1_uk_n1325 ) , .B1( u1_uk_n277 ) );
  NAND2_X1 u1_uk_U427 (.A1( u1_uk_K_r1_18 ) , .ZN( u1_uk_n1049 ) , .A2( u1_uk_n203 ) );
  BUF_X1 u1_uk_U43 (.Z( u1_uk_n220 ) , .A( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U434 (.ZN( u1_K5_16 ) , .B1( u1_uk_n129 ) , .A2( u1_uk_n1397 ) , .B2( u1_uk_n1410 ) , .A1( u1_uk_n251 ) );
  INV_X1 u1_uk_U436 (.ZN( u1_K2_28 ) , .A( u1_uk_n1028 ) );
  AOI22_X1 u1_uk_U437 (.B2( u1_uk_K_r0_15 ) , .A2( u1_uk_K_r0_49 ) , .ZN( u1_uk_n1028 ) , .A1( u1_uk_n164 ) , .B1( u1_uk_n220 ) );
  BUF_X1 u1_uk_U44 (.Z( u1_uk_n214 ) , .A( u1_uk_n286 ) );
  BUF_X1 u1_uk_U45 (.Z( u1_uk_n240 ) , .A( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U456 (.ZN( u1_K14_33 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1815 ) , .A2( u1_uk_n1833 ) , .A1( u1_uk_n251 ) );
  OAI22_X1 u1_uk_U459 (.ZN( u1_K7_33 ) , .A1( u1_uk_n141 ) , .B2( u1_uk_n1494 ) , .A2( u1_uk_n1514 ) , .B1( u1_uk_n279 ) );
  BUF_X1 u1_uk_U46 (.Z( u1_uk_n238 ) , .A( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U467 (.ZN( u1_K8_33 ) , .B2( u1_uk_n1528 ) , .A2( u1_uk_n1533 ) , .A1( u1_uk_n292 ) , .B1( u1_uk_n63 ) );
  BUF_X1 u1_uk_U47 (.Z( u1_uk_n217 ) , .A( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U471 (.ZN( u1_K13_37 ) , .B1( u1_uk_n100 ) , .B2( u1_uk_n1764 ) , .A2( u1_uk_n1776 ) , .A1( u1_uk_n271 ) );
  BUF_X1 u1_uk_U48 (.Z( u1_uk_n223 ) , .A( u1_uk_n277 ) );
  OAI21_X1 u1_uk_U483 (.ZN( u1_K14_29 ) , .B1( u1_uk_n155 ) , .B2( u1_uk_n1837 ) , .A( u1_uk_n954 ) );
  NAND2_X1 u1_uk_U484 (.A1( u1_uk_K_r12_44 ) , .A2( u1_uk_n164 ) , .ZN( u1_uk_n954 ) );
  OAI22_X1 u1_uk_U490 (.ZN( u1_K2_29 ) , .B1( u1_uk_n100 ) , .A2( u1_uk_n1267 ) , .B2( u1_uk_n1282 ) , .A1( u1_uk_n250 ) );
  OAI22_X1 u1_uk_U492 (.ZN( u1_K10_29 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1627 ) , .A2( u1_uk_n1655 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U493 (.ZN( u1_K9_29 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1595 ) , .A2( u1_uk_n1599 ) , .B1( u1_uk_n222 ) );
  INV_X1 u1_uk_U497 (.ZN( u1_K8_29 ) , .A( u1_uk_n1134 ) );
  AOI22_X1 u1_uk_U498 (.B2( u1_uk_K_r6_28 ) , .A2( u1_uk_K_r6_35 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1134 ) , .B1( u1_uk_n230 ) );
  INV_X1 u1_uk_U5 (.ZN( u1_uk_n163 ) , .A( u1_uk_n202 ) );
  BUF_X1 u1_uk_U50 (.Z( u1_uk_n191 ) , .A( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U507 (.ZN( u1_K3_2 ) , .B2( u1_uk_n1331 ) , .A2( u1_uk_n1336 ) , .A1( u1_uk_n208 ) , .B1( u1_uk_n94 ) );
  OAI21_X1 u1_uk_U511 (.ZN( u1_K7_2 ) , .A( u1_uk_n1116 ) , .B2( u1_uk_n1484 ) , .B1( u1_uk_n92 ) );
  NAND2_X1 u1_uk_U512 (.A1( u1_uk_K_r5_41 ) , .ZN( u1_uk_n1116 ) , .A2( u1_uk_n17 ) );
  OAI22_X1 u1_uk_U513 (.ZN( u1_K5_2 ) , .A1( u1_uk_n117 ) , .A2( u1_uk_n1397 ) , .B2( u1_uk_n1402 ) , .B1( u1_uk_n217 ) );
  OAI21_X1 u1_uk_U518 (.ZN( u1_K13_17 ) , .B1( u1_uk_n161 ) , .B2( u1_uk_n1773 ) , .A( u1_uk_n681 ) );
  NAND2_X1 u1_uk_U519 (.A1( u1_uk_K_r11_27 ) , .A2( u1_uk_n102 ) , .ZN( u1_uk_n681 ) );
  BUF_X1 u1_uk_U52 (.Z( u1_uk_n222 ) , .A( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U528 (.ZN( u1_K3_17 ) , .B2( u1_uk_n1317 ) , .A2( u1_uk_n1340 ) , .A1( u1_uk_n297 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U543 (.ZN( u1_K3_12 ) , .B2( u1_uk_n1336 ) , .A2( u1_uk_n1341 ) , .A1( u1_uk_n191 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U553 (.ZN( u1_K5_17 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1404 ) , .A2( u1_uk_n1424 ) , .B1( u1_uk_n277 ) );
  OAI22_X1 u1_uk_U557 (.ZN( u1_K14_36 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1800 ) , .A2( u1_uk_n1838 ) , .A1( u1_uk_n277 ) );
  INV_X1 u1_uk_U566 (.ZN( u1_K7_36 ) , .A( u1_uk_n1121 ) );
  AOI22_X1 u1_uk_U567 (.B2( u1_uk_K_r5_1 ) , .A2( u1_uk_K_r5_21 ) , .ZN( u1_uk_n1121 ) , .B1( u1_uk_n187 ) , .A1( u1_uk_n220 ) );
  BUF_X1 u1_uk_U57 (.Z( u1_uk_n286 ) , .A( u1_uk_n294 ) );
  OAI22_X1 u1_uk_U576 (.ZN( u1_K8_36 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1554 ) , .A2( u1_uk_n1560 ) , .A1( u1_uk_n217 ) );
  BUF_X1 u1_uk_U59 (.Z( u1_uk_n279 ) , .A( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U598 (.ZN( u1_K3_22 ) , .B2( u1_uk_n1311 ) , .A2( u1_uk_n1346 ) , .A1( u1_uk_n147 ) , .B1( u1_uk_n191 ) );
  BUF_X1 u1_uk_U60 (.Z( u1_uk_n271 ) , .A( u1_uk_n297 ) );
  BUF_X1 u1_uk_U61 (.Z( u1_uk_n277 ) , .A( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U614 (.ZN( u1_K8_35 ) , .B2( u1_uk_n1541 ) , .A2( u1_uk_n1547 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n99 ) );
  OAI21_X1 u1_uk_U615 (.ZN( u1_K7_35 ) , .A( u1_uk_n1120 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1482 ) );
  NAND2_X1 u1_uk_U616 (.A1( u1_uk_K_r5_37 ) , .ZN( u1_uk_n1120 ) , .A2( u1_uk_n17 ) );
  BUF_X1 u1_uk_U62 (.Z( u1_uk_n292 ) , .A( u1_uk_n294 ) );
  INV_X1 u1_uk_U620 (.ZN( u1_K14_35 ) , .A( u1_uk_n956 ) );
  AOI22_X1 u1_uk_U621 (.B2( u1_uk_K_r12_1 ) , .A2( u1_uk_K_r12_7 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n242 ) , .ZN( u1_uk_n956 ) );
  OAI22_X1 u1_uk_U639 (.ZN( u1_K3_11 ) , .A2( u1_uk_n1310 ) , .B2( u1_uk_n1315 ) , .A1( u1_uk_n146 ) , .B1( u1_uk_n191 ) );
  OAI22_X1 u1_uk_U664 (.ZN( u1_K9_25 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1608 ) , .A2( u1_uk_n1615 ) , .B1( u1_uk_n292 ) );
  OAI21_X1 u1_uk_U671 (.ZN( u1_K13_43 ) , .B2( u1_uk_n1792 ) , .B1( u1_uk_n191 ) , .A( u1_uk_n946 ) );
  NAND2_X1 u1_uk_U672 (.A1( u1_uk_K_r11_29 ) , .A2( u1_uk_n294 ) , .ZN( u1_uk_n946 ) );
  OAI21_X1 u1_uk_U692 (.ZN( u1_K2_25 ) , .A( u1_uk_n1026 ) , .B2( u1_uk_n1294 ) , .B1( u1_uk_n162 ) );
  NAND2_X1 u1_uk_U693 (.A1( u1_uk_K_r0_22 ) , .ZN( u1_uk_n1026 ) , .A2( u1_uk_n109 ) );
  OAI22_X1 u1_uk_U696 (.ZN( u1_K10_25 ) , .A1( u1_uk_n109 ) , .A2( u1_uk_n1623 ) , .B2( u1_uk_n1641 ) , .B1( u1_uk_n291 ) );
  OAI22_X1 u1_uk_U697 (.ZN( u1_K8_25 ) , .B1( u1_uk_n102 ) , .B2( u1_uk_n1563 ) , .A2( u1_uk_n1568 ) , .A1( u1_uk_n214 ) );
  INV_X1 u1_uk_U71 (.ZN( u1_K8_34 ) , .A( u1_uk_n1137 ) );
  AOI22_X1 u1_uk_U72 (.B2( u1_uk_K_r6_14 ) , .A2( u1_uk_K_r6_21 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1137 ) , .B1( u1_uk_n214 ) );
  OAI22_X1 u1_uk_U724 (.ZN( u1_K8_32 ) , .B2( u1_uk_n1556 ) , .A2( u1_uk_n1563 ) , .A1( u1_uk_n271 ) , .B1( u1_uk_n93 ) );
  INV_X1 u1_uk_U73 (.ZN( u1_K7_34 ) , .A( u1_uk_n1119 ) );
  OAI22_X1 u1_uk_U730 (.ZN( u1_K14_32 ) , .B1( u1_uk_n109 ) , .B2( u1_uk_n1799 ) , .A2( u1_uk_n1837 ) , .A1( u1_uk_n286 ) );
  OAI22_X1 u1_uk_U734 (.ZN( u1_K13_42 ) , .A1( u1_uk_n145 ) , .B2( u1_uk_n1763 ) , .A2( u1_uk_n1769 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U739 (.ZN( u1_K2_42 ) , .B2( u1_uk_n1296 ) , .A2( u1_uk_n1304 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n93 ) );
  AOI22_X1 u1_uk_U74 (.B2( u1_uk_K_r5_0 ) , .A2( u1_uk_K_r5_35 ) , .A1( u1_uk_n110 ) , .ZN( u1_uk_n1119 ) , .B1( u1_uk_n209 ) );
  OAI21_X1 u1_uk_U748 (.ZN( u1_K14_27 ) , .B2( u1_uk_n1839 ) , .B1( u1_uk_n63 ) , .A( u1_uk_n953 ) );
  NAND2_X1 u1_uk_U749 (.A1( u1_uk_K_r12_42 ) , .A2( u1_uk_n10 ) , .ZN( u1_uk_n953 ) );
  OAI21_X1 u1_uk_U751 (.ZN( u1_K10_27 ) , .B1( u1_uk_n11 ) , .B2( u1_uk_n1632 ) , .A( u1_uk_n335 ) );
  NAND2_X1 u1_uk_U752 (.A1( u1_uk_K_r8_43 ) , .A2( u1_uk_n27 ) , .ZN( u1_uk_n335 ) );
  OAI22_X1 u1_uk_U753 (.ZN( u1_K8_27 ) , .B1( u1_uk_n148 ) , .B2( u1_uk_n1529 ) , .A2( u1_uk_n1534 ) , .A1( u1_uk_n202 ) );
  INV_X1 u1_uk_U76 (.ZN( u1_K14_34 ) , .A( u1_uk_n955 ) );
  AOI22_X1 u1_uk_U77 (.B2( u1_uk_K_r12_30 ) , .A2( u1_uk_K_r12_36 ) , .B1( u1_uk_n163 ) , .A1( u1_uk_n279 ) , .ZN( u1_uk_n955 ) );
  INV_X1 u1_uk_U781 (.ZN( u1_K13_13 ) , .A( u1_uk_n677 ) );
  AOI22_X1 u1_uk_U782 (.B2( u1_uk_K_r11_11 ) , .A2( u1_uk_K_r11_6 ) , .A1( u1_uk_n109 ) , .B1( u1_uk_n240 ) , .ZN( u1_uk_n677 ) );
  INV_X1 u1_uk_U792 (.ZN( u1_K2_27 ) , .A( u1_uk_n1027 ) );
  AOI22_X1 u1_uk_U793 (.B2( u1_uk_K_r0_28 ) , .A2( u1_uk_K_r0_7 ) , .ZN( u1_uk_n1027 ) , .A1( u1_uk_n129 ) , .B1( u1_uk_n252 ) );
  INV_X1 u1_uk_U800 (.ZN( u1_K9_27 ) , .A( u1_uk_n1159 ) );
  AOI22_X1 u1_uk_U801 (.B2( u1_uk_K_r7_2 ) , .A2( u1_uk_K_r7_9 ) , .B1( u1_uk_n100 ) , .ZN( u1_uk_n1159 ) , .A1( u1_uk_n279 ) );
  OAI22_X1 u1_uk_U812 (.ZN( u1_K5_18 ) , .A2( u1_uk_n1399 ) , .B2( u1_uk_n1436 ) , .B1( u1_uk_n146 ) , .A1( u1_uk_n188 ) );
  OAI21_X1 u1_uk_U815 (.ZN( u1_K13_18 ) , .B2( u1_uk_n1780 ) , .B1( u1_uk_n231 ) , .A( u1_uk_n682 ) );
  NAND2_X1 u1_uk_U816 (.A1( u1_uk_K_r11_20 ) , .A2( u1_uk_n291 ) , .ZN( u1_uk_n682 ) );
  OAI22_X1 u1_uk_U825 (.ZN( u1_K3_20 ) , .B2( u1_uk_n1320 ) , .A2( u1_uk_n1326 ) , .A1( u1_uk_n242 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U849 (.ZN( u1_K7_3 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1495 ) , .A2( u1_uk_n1517 ) , .B1( u1_uk_n217 ) );
  INV_X1 u1_uk_U851 (.ZN( u1_K7_6 ) , .A( u1_uk_n1125 ) );
  AOI22_X1 u1_uk_U852 (.B2( u1_uk_K_r5_39 ) , .A2( u1_uk_K_r5_4 ) , .ZN( u1_uk_n1125 ) , .B1( u1_uk_n182 ) , .A1( u1_uk_n188 ) );
  OAI21_X1 u1_uk_U855 (.ZN( u1_K3_3 ) , .A( u1_uk_n1043 ) , .B2( u1_uk_n1348 ) , .B1( u1_uk_n242 ) );
  NAND2_X1 u1_uk_U856 (.A1( u1_uk_K_r1_47 ) , .ZN( u1_uk_n1043 ) , .A2( u1_uk_n292 ) );
  OAI22_X1 u1_uk_U866 (.ZN( u1_K3_18 ) , .B2( u1_uk_n1325 ) , .A2( u1_uk_n1332 ) , .A1( u1_uk_n240 ) , .B1( u1_uk_n31 ) );
  OAI22_X1 u1_uk_U884 (.ZN( u1_K3_10 ) , .B2( u1_uk_n1316 ) , .A2( u1_uk_n1321 ) , .A1( u1_uk_n217 ) , .B1( u1_uk_n63 ) );
  OAI22_X1 u1_uk_U886 (.ZN( u1_K13_45 ) , .B1( u1_uk_n162 ) , .B2( u1_uk_n1755 ) , .A2( u1_uk_n1793 ) , .A1( u1_uk_n271 ) );
  OAI22_X1 u1_uk_U896 (.ZN( u1_K5_3 ) , .B2( u1_uk_n1404 ) , .A2( u1_uk_n1411 ) , .A1( u1_uk_n230 ) , .B1( u1_uk_n93 ) );
  OAI22_X1 u1_uk_U902 (.ZN( u1_K3_21 ) , .B2( u1_uk_n1321 ) , .A2( u1_uk_n1346 ) , .A1( u1_uk_n250 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U911 (.ZN( u1_K5_13 ) , .B1( u1_uk_n117 ) , .B2( u1_uk_n1405 ) , .A2( u1_uk_n1436 ) , .A1( u1_uk_n297 ) );
  OAI22_X1 u1_uk_U912 (.ZN( u1_K5_14 ) , .B2( u1_uk_n1403 ) , .B1( u1_uk_n141 ) , .A2( u1_uk_n1410 ) , .A1( u1_uk_n220 ) );
  OAI22_X1 u1_uk_U914 (.ZN( u1_K3_13 ) , .B2( u1_uk_n1319 ) , .A2( u1_uk_n1324 ) , .A1( u1_uk_n298 ) , .B1( u1_uk_n60 ) );
  OAI22_X1 u1_uk_U927 (.ZN( u1_K2_39 ) , .A2( u1_uk_n1266 ) , .B2( u1_uk_n1281 ) , .A1( u1_uk_n222 ) , .B1( u1_uk_n99 ) );
  OAI22_X1 u1_uk_U93 (.ZN( u1_K3_23 ) , .A1( u1_uk_n118 ) , .A2( u1_uk_n1311 ) , .B2( u1_uk_n1316 ) , .B1( u1_uk_n202 ) );
  OAI22_X1 u1_uk_U967 (.ZN( u1_K13_38 ) , .A1( u1_uk_n146 ) , .B2( u1_uk_n1785 ) , .A2( u1_uk_n1791 ) , .B1( u1_uk_n231 ) );
  OAI22_X1 u1_uk_U968 (.ZN( u1_K2_38 ) , .A1( u1_uk_n110 ) , .B2( u1_uk_n1276 ) , .A2( u1_uk_n1295 ) , .B1( u1_uk_n238 ) );
  OAI22_X1 u1_uk_U970 (.ZN( u1_K2_37 ) , .A2( u1_uk_n1267 ) , .B2( u1_uk_n1294 ) , .B1( u1_uk_n252 ) , .A1( u1_uk_n83 ) );
  OAI22_X1 u1_uk_U982 (.ZN( u1_K3_6 ) , .A2( u1_uk_n1312 ) , .B2( u1_uk_n1317 ) , .A1( u1_uk_n182 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U985 (.ZN( u1_K3_7 ) , .A1( u1_uk_n118 ) , .B2( u1_uk_n1323 ) , .A2( u1_uk_n1341 ) , .B1( u1_uk_n208 ) );
  OAI22_X1 u1_uk_U989 (.ZN( u1_K14_25 ) , .A1( u1_uk_n142 ) , .B2( u1_uk_n1800 ) , .A2( u1_uk_n1806 ) , .B1( u1_uk_n222 ) );
  INV_X1 u1_uk_U99 (.ZN( u1_K2_41 ) , .A( u1_uk_n1031 ) );
  XOR2_X1 u2_U350 (.B( u2_L5_26 ) , .Z( u2_N217 ) , .A( u2_out6_26 ) );
  XOR2_X1 u2_U356 (.B( u2_L5_20 ) , .Z( u2_N211 ) , .A( u2_out6_20 ) );
  XOR2_X1 u2_U367 (.B( u2_L5_10 ) , .Z( u2_N201 ) , .A( u2_out6_10 ) );
  XOR2_X1 u2_U378 (.B( u2_L5_1 ) , .Z( u2_N192 ) , .A( u2_out6_1 ) );
  XOR2_X1 u2_U487 (.Z( u2_FP_5 ) , .B( u2_L14_5 ) , .A( u2_out15_5 ) );
  XOR2_X1 u2_U496 (.Z( u2_FP_27 ) , .B( u2_L14_27 ) , .A( u2_out15_27 ) );
  XOR2_X1 u2_U502 (.Z( u2_FP_21 ) , .B( u2_L14_21 ) , .A( u2_out15_21 ) );
  XOR2_X1 u2_U509 (.Z( u2_FP_15 ) , .B( u2_L14_15 ) , .A( u2_out15_15 ) );
  XOR2_X1 u2_u15_U10 (.A( u2_FP_62 ) , .B( u2_K16_45 ) , .Z( u2_u15_X_45 ) );
  XOR2_X1 u2_u15_U11 (.A( u2_FP_61 ) , .B( u2_K16_44 ) , .Z( u2_u15_X_44 ) );
  XOR2_X1 u2_u15_U12 (.A( u2_FP_60 ) , .B( u2_K16_43 ) , .Z( u2_u15_X_43 ) );
  XOR2_X1 u2_u15_U7 (.A( u2_FP_33 ) , .B( u2_K16_48 ) , .Z( u2_u15_X_48 ) );
  XOR2_X1 u2_u15_U8 (.A( u2_FP_64 ) , .B( u2_K16_47 ) , .Z( u2_u15_X_47 ) );
  XOR2_X1 u2_u15_U9 (.A( u2_FP_63 ) , .B( u2_K16_46 ) , .Z( u2_u15_X_46 ) );
  OAI21_X1 u2_u15_u7_U10 (.A( u2_u15_u7_n161 ) , .B1( u2_u15_u7_n168 ) , .B2( u2_u15_u7_n173 ) , .ZN( u2_u15_u7_n91 ) );
  AOI211_X1 u2_u15_u7_U11 (.A( u2_u15_u7_n117 ) , .ZN( u2_u15_u7_n118 ) , .C2( u2_u15_u7_n126 ) , .C1( u2_u15_u7_n177 ) , .B( u2_u15_u7_n180 ) );
  OAI22_X1 u2_u15_u7_U12 (.B1( u2_u15_u7_n115 ) , .ZN( u2_u15_u7_n117 ) , .A2( u2_u15_u7_n133 ) , .A1( u2_u15_u7_n137 ) , .B2( u2_u15_u7_n162 ) );
  INV_X1 u2_u15_u7_U13 (.A( u2_u15_u7_n116 ) , .ZN( u2_u15_u7_n180 ) );
  NOR3_X1 u2_u15_u7_U14 (.ZN( u2_u15_u7_n115 ) , .A3( u2_u15_u7_n145 ) , .A2( u2_u15_u7_n168 ) , .A1( u2_u15_u7_n169 ) );
  OAI211_X1 u2_u15_u7_U15 (.B( u2_u15_u7_n122 ) , .A( u2_u15_u7_n123 ) , .C2( u2_u15_u7_n124 ) , .ZN( u2_u15_u7_n154 ) , .C1( u2_u15_u7_n162 ) );
  AOI222_X1 u2_u15_u7_U16 (.ZN( u2_u15_u7_n122 ) , .C2( u2_u15_u7_n126 ) , .C1( u2_u15_u7_n145 ) , .B1( u2_u15_u7_n161 ) , .A2( u2_u15_u7_n165 ) , .B2( u2_u15_u7_n170 ) , .A1( u2_u15_u7_n176 ) );
  INV_X1 u2_u15_u7_U17 (.A( u2_u15_u7_n133 ) , .ZN( u2_u15_u7_n176 ) );
  NOR3_X1 u2_u15_u7_U18 (.A2( u2_u15_u7_n134 ) , .A1( u2_u15_u7_n135 ) , .ZN( u2_u15_u7_n136 ) , .A3( u2_u15_u7_n171 ) );
  NOR2_X1 u2_u15_u7_U19 (.A1( u2_u15_u7_n130 ) , .A2( u2_u15_u7_n134 ) , .ZN( u2_u15_u7_n153 ) );
  INV_X1 u2_u15_u7_U20 (.A( u2_u15_u7_n101 ) , .ZN( u2_u15_u7_n165 ) );
  NOR2_X1 u2_u15_u7_U21 (.ZN( u2_u15_u7_n111 ) , .A2( u2_u15_u7_n134 ) , .A1( u2_u15_u7_n169 ) );
  AOI21_X1 u2_u15_u7_U22 (.ZN( u2_u15_u7_n104 ) , .B2( u2_u15_u7_n112 ) , .B1( u2_u15_u7_n127 ) , .A( u2_u15_u7_n164 ) );
  AOI21_X1 u2_u15_u7_U23 (.ZN( u2_u15_u7_n106 ) , .B1( u2_u15_u7_n133 ) , .B2( u2_u15_u7_n146 ) , .A( u2_u15_u7_n162 ) );
  AOI21_X1 u2_u15_u7_U24 (.A( u2_u15_u7_n101 ) , .ZN( u2_u15_u7_n107 ) , .B2( u2_u15_u7_n128 ) , .B1( u2_u15_u7_n175 ) );
  INV_X1 u2_u15_u7_U25 (.A( u2_u15_u7_n138 ) , .ZN( u2_u15_u7_n171 ) );
  INV_X1 u2_u15_u7_U26 (.A( u2_u15_u7_n131 ) , .ZN( u2_u15_u7_n177 ) );
  INV_X1 u2_u15_u7_U27 (.A( u2_u15_u7_n110 ) , .ZN( u2_u15_u7_n174 ) );
  NAND2_X1 u2_u15_u7_U28 (.A1( u2_u15_u7_n129 ) , .A2( u2_u15_u7_n132 ) , .ZN( u2_u15_u7_n149 ) );
  NAND2_X1 u2_u15_u7_U29 (.A1( u2_u15_u7_n113 ) , .A2( u2_u15_u7_n124 ) , .ZN( u2_u15_u7_n130 ) );
  INV_X1 u2_u15_u7_U3 (.A( u2_u15_u7_n111 ) , .ZN( u2_u15_u7_n170 ) );
  INV_X1 u2_u15_u7_U30 (.A( u2_u15_u7_n112 ) , .ZN( u2_u15_u7_n173 ) );
  INV_X1 u2_u15_u7_U31 (.A( u2_u15_u7_n128 ) , .ZN( u2_u15_u7_n168 ) );
  INV_X1 u2_u15_u7_U32 (.A( u2_u15_u7_n148 ) , .ZN( u2_u15_u7_n169 ) );
  INV_X1 u2_u15_u7_U33 (.A( u2_u15_u7_n127 ) , .ZN( u2_u15_u7_n179 ) );
  NOR2_X1 u2_u15_u7_U34 (.ZN( u2_u15_u7_n101 ) , .A2( u2_u15_u7_n150 ) , .A1( u2_u15_u7_n156 ) );
  AOI211_X1 u2_u15_u7_U35 (.B( u2_u15_u7_n154 ) , .A( u2_u15_u7_n155 ) , .C1( u2_u15_u7_n156 ) , .ZN( u2_u15_u7_n157 ) , .C2( u2_u15_u7_n172 ) );
  INV_X1 u2_u15_u7_U36 (.A( u2_u15_u7_n153 ) , .ZN( u2_u15_u7_n172 ) );
  AOI211_X1 u2_u15_u7_U37 (.B( u2_u15_u7_n139 ) , .A( u2_u15_u7_n140 ) , .C2( u2_u15_u7_n141 ) , .ZN( u2_u15_u7_n142 ) , .C1( u2_u15_u7_n156 ) );
  NAND4_X1 u2_u15_u7_U38 (.A3( u2_u15_u7_n127 ) , .A2( u2_u15_u7_n128 ) , .A1( u2_u15_u7_n129 ) , .ZN( u2_u15_u7_n141 ) , .A4( u2_u15_u7_n147 ) );
  AOI21_X1 u2_u15_u7_U39 (.A( u2_u15_u7_n137 ) , .B1( u2_u15_u7_n138 ) , .ZN( u2_u15_u7_n139 ) , .B2( u2_u15_u7_n146 ) );
  INV_X1 u2_u15_u7_U4 (.A( u2_u15_u7_n149 ) , .ZN( u2_u15_u7_n175 ) );
  OAI22_X1 u2_u15_u7_U40 (.B1( u2_u15_u7_n136 ) , .ZN( u2_u15_u7_n140 ) , .A1( u2_u15_u7_n153 ) , .B2( u2_u15_u7_n162 ) , .A2( u2_u15_u7_n164 ) );
  AOI21_X1 u2_u15_u7_U41 (.ZN( u2_u15_u7_n123 ) , .B1( u2_u15_u7_n165 ) , .B2( u2_u15_u7_n177 ) , .A( u2_u15_u7_n97 ) );
  AOI21_X1 u2_u15_u7_U42 (.B2( u2_u15_u7_n113 ) , .B1( u2_u15_u7_n124 ) , .A( u2_u15_u7_n125 ) , .ZN( u2_u15_u7_n97 ) );
  INV_X1 u2_u15_u7_U43 (.A( u2_u15_u7_n125 ) , .ZN( u2_u15_u7_n161 ) );
  INV_X1 u2_u15_u7_U44 (.A( u2_u15_u7_n152 ) , .ZN( u2_u15_u7_n162 ) );
  AOI22_X1 u2_u15_u7_U45 (.A2( u2_u15_u7_n114 ) , .ZN( u2_u15_u7_n119 ) , .B1( u2_u15_u7_n130 ) , .A1( u2_u15_u7_n156 ) , .B2( u2_u15_u7_n165 ) );
  NAND2_X1 u2_u15_u7_U46 (.A2( u2_u15_u7_n112 ) , .ZN( u2_u15_u7_n114 ) , .A1( u2_u15_u7_n175 ) );
  AOI22_X1 u2_u15_u7_U47 (.B2( u2_u15_u7_n149 ) , .B1( u2_u15_u7_n150 ) , .A2( u2_u15_u7_n151 ) , .A1( u2_u15_u7_n152 ) , .ZN( u2_u15_u7_n158 ) );
  AND2_X1 u2_u15_u7_U48 (.ZN( u2_u15_u7_n145 ) , .A2( u2_u15_u7_n98 ) , .A1( u2_u15_u7_n99 ) );
  NOR2_X1 u2_u15_u7_U49 (.ZN( u2_u15_u7_n137 ) , .A1( u2_u15_u7_n150 ) , .A2( u2_u15_u7_n161 ) );
  INV_X1 u2_u15_u7_U5 (.A( u2_u15_u7_n154 ) , .ZN( u2_u15_u7_n178 ) );
  AOI21_X1 u2_u15_u7_U50 (.ZN( u2_u15_u7_n105 ) , .B2( u2_u15_u7_n110 ) , .A( u2_u15_u7_n125 ) , .B1( u2_u15_u7_n147 ) );
  NAND2_X1 u2_u15_u7_U51 (.ZN( u2_u15_u7_n146 ) , .A1( u2_u15_u7_n95 ) , .A2( u2_u15_u7_n98 ) );
  NAND2_X1 u2_u15_u7_U52 (.A2( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n147 ) , .A1( u2_u15_u7_n93 ) );
  NAND2_X1 u2_u15_u7_U53 (.A1( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n127 ) , .A2( u2_u15_u7_n99 ) );
  OR2_X1 u2_u15_u7_U54 (.ZN( u2_u15_u7_n126 ) , .A2( u2_u15_u7_n152 ) , .A1( u2_u15_u7_n156 ) );
  NAND2_X1 u2_u15_u7_U55 (.A2( u2_u15_u7_n102 ) , .A1( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n133 ) );
  NAND2_X1 u2_u15_u7_U56 (.ZN( u2_u15_u7_n112 ) , .A2( u2_u15_u7_n96 ) , .A1( u2_u15_u7_n99 ) );
  NAND2_X1 u2_u15_u7_U57 (.A2( u2_u15_u7_n102 ) , .ZN( u2_u15_u7_n128 ) , .A1( u2_u15_u7_n98 ) );
  NAND2_X1 u2_u15_u7_U58 (.A1( u2_u15_u7_n100 ) , .ZN( u2_u15_u7_n113 ) , .A2( u2_u15_u7_n93 ) );
  NAND2_X1 u2_u15_u7_U59 (.A2( u2_u15_u7_n102 ) , .ZN( u2_u15_u7_n124 ) , .A1( u2_u15_u7_n96 ) );
  AOI211_X1 u2_u15_u7_U6 (.ZN( u2_u15_u7_n116 ) , .A( u2_u15_u7_n155 ) , .C1( u2_u15_u7_n161 ) , .C2( u2_u15_u7_n171 ) , .B( u2_u15_u7_n94 ) );
  NAND2_X1 u2_u15_u7_U60 (.ZN( u2_u15_u7_n110 ) , .A1( u2_u15_u7_n95 ) , .A2( u2_u15_u7_n96 ) );
  INV_X1 u2_u15_u7_U61 (.A( u2_u15_u7_n150 ) , .ZN( u2_u15_u7_n164 ) );
  AND2_X1 u2_u15_u7_U62 (.ZN( u2_u15_u7_n134 ) , .A1( u2_u15_u7_n93 ) , .A2( u2_u15_u7_n98 ) );
  NAND2_X1 u2_u15_u7_U63 (.A1( u2_u15_u7_n100 ) , .A2( u2_u15_u7_n102 ) , .ZN( u2_u15_u7_n129 ) );
  NAND2_X1 u2_u15_u7_U64 (.A2( u2_u15_u7_n103 ) , .ZN( u2_u15_u7_n131 ) , .A1( u2_u15_u7_n95 ) );
  NAND2_X1 u2_u15_u7_U65 (.A1( u2_u15_u7_n100 ) , .ZN( u2_u15_u7_n138 ) , .A2( u2_u15_u7_n99 ) );
  NAND2_X1 u2_u15_u7_U66 (.ZN( u2_u15_u7_n132 ) , .A1( u2_u15_u7_n93 ) , .A2( u2_u15_u7_n96 ) );
  NAND2_X1 u2_u15_u7_U67 (.A1( u2_u15_u7_n100 ) , .ZN( u2_u15_u7_n148 ) , .A2( u2_u15_u7_n95 ) );
  NOR2_X1 u2_u15_u7_U68 (.A2( u2_u15_X_47 ) , .ZN( u2_u15_u7_n150 ) , .A1( u2_u15_u7_n163 ) );
  NOR2_X1 u2_u15_u7_U69 (.A2( u2_u15_X_43 ) , .A1( u2_u15_X_44 ) , .ZN( u2_u15_u7_n103 ) );
  OAI222_X1 u2_u15_u7_U7 (.C2( u2_u15_u7_n101 ) , .B2( u2_u15_u7_n111 ) , .A1( u2_u15_u7_n113 ) , .C1( u2_u15_u7_n146 ) , .A2( u2_u15_u7_n162 ) , .B1( u2_u15_u7_n164 ) , .ZN( u2_u15_u7_n94 ) );
  NOR2_X1 u2_u15_u7_U70 (.A2( u2_u15_X_48 ) , .A1( u2_u15_u7_n166 ) , .ZN( u2_u15_u7_n95 ) );
  NOR2_X1 u2_u15_u7_U71 (.A2( u2_u15_X_45 ) , .A1( u2_u15_X_48 ) , .ZN( u2_u15_u7_n99 ) );
  NOR2_X1 u2_u15_u7_U72 (.A2( u2_u15_X_44 ) , .A1( u2_u15_u7_n167 ) , .ZN( u2_u15_u7_n98 ) );
  NOR2_X1 u2_u15_u7_U73 (.A2( u2_u15_X_46 ) , .A1( u2_u15_X_47 ) , .ZN( u2_u15_u7_n152 ) );
  AND2_X1 u2_u15_u7_U74 (.A1( u2_u15_X_47 ) , .ZN( u2_u15_u7_n156 ) , .A2( u2_u15_u7_n163 ) );
  NAND2_X1 u2_u15_u7_U75 (.A2( u2_u15_X_46 ) , .A1( u2_u15_X_47 ) , .ZN( u2_u15_u7_n125 ) );
  AND2_X1 u2_u15_u7_U76 (.A2( u2_u15_X_45 ) , .A1( u2_u15_X_48 ) , .ZN( u2_u15_u7_n102 ) );
  AND2_X1 u2_u15_u7_U77 (.A2( u2_u15_X_43 ) , .A1( u2_u15_X_44 ) , .ZN( u2_u15_u7_n96 ) );
  AND2_X1 u2_u15_u7_U78 (.A1( u2_u15_X_44 ) , .ZN( u2_u15_u7_n100 ) , .A2( u2_u15_u7_n167 ) );
  AND2_X1 u2_u15_u7_U79 (.A1( u2_u15_X_48 ) , .A2( u2_u15_u7_n166 ) , .ZN( u2_u15_u7_n93 ) );
  OAI221_X1 u2_u15_u7_U8 (.C1( u2_u15_u7_n101 ) , .C2( u2_u15_u7_n147 ) , .ZN( u2_u15_u7_n155 ) , .B2( u2_u15_u7_n162 ) , .A( u2_u15_u7_n91 ) , .B1( u2_u15_u7_n92 ) );
  INV_X1 u2_u15_u7_U80 (.A( u2_u15_X_46 ) , .ZN( u2_u15_u7_n163 ) );
  INV_X1 u2_u15_u7_U81 (.A( u2_u15_X_45 ) , .ZN( u2_u15_u7_n166 ) );
  INV_X1 u2_u15_u7_U82 (.A( u2_u15_X_43 ) , .ZN( u2_u15_u7_n167 ) );
  NAND4_X1 u2_u15_u7_U83 (.ZN( u2_out15_5 ) , .A4( u2_u15_u7_n108 ) , .A3( u2_u15_u7_n109 ) , .A1( u2_u15_u7_n116 ) , .A2( u2_u15_u7_n123 ) );
  AOI22_X1 u2_u15_u7_U84 (.ZN( u2_u15_u7_n109 ) , .A2( u2_u15_u7_n126 ) , .B2( u2_u15_u7_n145 ) , .B1( u2_u15_u7_n156 ) , .A1( u2_u15_u7_n171 ) );
  NOR4_X1 u2_u15_u7_U85 (.A4( u2_u15_u7_n104 ) , .A3( u2_u15_u7_n105 ) , .A2( u2_u15_u7_n106 ) , .A1( u2_u15_u7_n107 ) , .ZN( u2_u15_u7_n108 ) );
  NAND4_X1 u2_u15_u7_U86 (.ZN( u2_out15_27 ) , .A4( u2_u15_u7_n118 ) , .A3( u2_u15_u7_n119 ) , .A2( u2_u15_u7_n120 ) , .A1( u2_u15_u7_n121 ) );
  OAI21_X1 u2_u15_u7_U87 (.ZN( u2_u15_u7_n121 ) , .B2( u2_u15_u7_n145 ) , .A( u2_u15_u7_n150 ) , .B1( u2_u15_u7_n174 ) );
  OAI21_X1 u2_u15_u7_U88 (.ZN( u2_u15_u7_n120 ) , .A( u2_u15_u7_n161 ) , .B2( u2_u15_u7_n170 ) , .B1( u2_u15_u7_n179 ) );
  NAND4_X1 u2_u15_u7_U89 (.ZN( u2_out15_21 ) , .A4( u2_u15_u7_n157 ) , .A3( u2_u15_u7_n158 ) , .A2( u2_u15_u7_n159 ) , .A1( u2_u15_u7_n160 ) );
  AND3_X1 u2_u15_u7_U9 (.A3( u2_u15_u7_n110 ) , .A2( u2_u15_u7_n127 ) , .A1( u2_u15_u7_n132 ) , .ZN( u2_u15_u7_n92 ) );
  OAI21_X1 u2_u15_u7_U90 (.B1( u2_u15_u7_n145 ) , .ZN( u2_u15_u7_n160 ) , .A( u2_u15_u7_n161 ) , .B2( u2_u15_u7_n177 ) );
  OAI21_X1 u2_u15_u7_U91 (.ZN( u2_u15_u7_n159 ) , .A( u2_u15_u7_n165 ) , .B2( u2_u15_u7_n171 ) , .B1( u2_u15_u7_n174 ) );
  NAND4_X1 u2_u15_u7_U92 (.ZN( u2_out15_15 ) , .A4( u2_u15_u7_n142 ) , .A3( u2_u15_u7_n143 ) , .A2( u2_u15_u7_n144 ) , .A1( u2_u15_u7_n178 ) );
  OR2_X1 u2_u15_u7_U93 (.A2( u2_u15_u7_n125 ) , .A1( u2_u15_u7_n129 ) , .ZN( u2_u15_u7_n144 ) );
  AOI22_X1 u2_u15_u7_U94 (.A2( u2_u15_u7_n126 ) , .ZN( u2_u15_u7_n143 ) , .B2( u2_u15_u7_n165 ) , .B1( u2_u15_u7_n173 ) , .A1( u2_u15_u7_n174 ) );
  NAND3_X1 u2_u15_u7_U95 (.A3( u2_u15_u7_n146 ) , .A2( u2_u15_u7_n147 ) , .A1( u2_u15_u7_n148 ) , .ZN( u2_u15_u7_n151 ) );
  NAND3_X1 u2_u15_u7_U96 (.A3( u2_u15_u7_n131 ) , .A2( u2_u15_u7_n132 ) , .A1( u2_u15_u7_n133 ) , .ZN( u2_u15_u7_n135 ) );
  XOR2_X1 u2_u6_U33 (.B( u2_K7_24 ) , .A( u2_R5_17 ) , .Z( u2_u6_X_24 ) );
  XOR2_X1 u2_u6_U34 (.B( u2_K7_23 ) , .A( u2_R5_16 ) , .Z( u2_u6_X_23 ) );
  XOR2_X1 u2_u6_U35 (.B( u2_K7_22 ) , .A( u2_R5_15 ) , .Z( u2_u6_X_22 ) );
  XOR2_X1 u2_u6_U36 (.B( u2_K7_21 ) , .A( u2_R5_14 ) , .Z( u2_u6_X_21 ) );
  XOR2_X1 u2_u6_U37 (.B( u2_K7_20 ) , .A( u2_R5_13 ) , .Z( u2_u6_X_20 ) );
  XOR2_X1 u2_u6_U39 (.B( u2_K7_19 ) , .A( u2_R5_12 ) , .Z( u2_u6_X_19 ) );
  OAI22_X1 u2_u6_u3_U10 (.B1( u2_u6_u3_n113 ) , .A2( u2_u6_u3_n135 ) , .A1( u2_u6_u3_n150 ) , .B2( u2_u6_u3_n164 ) , .ZN( u2_u6_u3_n98 ) );
  OAI211_X1 u2_u6_u3_U11 (.B( u2_u6_u3_n106 ) , .ZN( u2_u6_u3_n119 ) , .C2( u2_u6_u3_n128 ) , .C1( u2_u6_u3_n167 ) , .A( u2_u6_u3_n181 ) );
  AOI221_X1 u2_u6_u3_U12 (.C1( u2_u6_u3_n105 ) , .ZN( u2_u6_u3_n106 ) , .A( u2_u6_u3_n131 ) , .B2( u2_u6_u3_n132 ) , .C2( u2_u6_u3_n133 ) , .B1( u2_u6_u3_n169 ) );
  INV_X1 u2_u6_u3_U13 (.ZN( u2_u6_u3_n181 ) , .A( u2_u6_u3_n98 ) );
  NAND2_X1 u2_u6_u3_U14 (.ZN( u2_u6_u3_n105 ) , .A2( u2_u6_u3_n130 ) , .A1( u2_u6_u3_n155 ) );
  NOR2_X1 u2_u6_u3_U15 (.ZN( u2_u6_u3_n126 ) , .A2( u2_u6_u3_n150 ) , .A1( u2_u6_u3_n164 ) );
  AOI21_X1 u2_u6_u3_U16 (.ZN( u2_u6_u3_n112 ) , .B2( u2_u6_u3_n146 ) , .B1( u2_u6_u3_n155 ) , .A( u2_u6_u3_n167 ) );
  NAND2_X1 u2_u6_u3_U17 (.A1( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n142 ) , .A2( u2_u6_u3_n164 ) );
  NAND2_X1 u2_u6_u3_U18 (.ZN( u2_u6_u3_n132 ) , .A2( u2_u6_u3_n152 ) , .A1( u2_u6_u3_n156 ) );
  AND2_X1 u2_u6_u3_U19 (.A2( u2_u6_u3_n113 ) , .A1( u2_u6_u3_n114 ) , .ZN( u2_u6_u3_n151 ) );
  INV_X1 u2_u6_u3_U20 (.A( u2_u6_u3_n133 ) , .ZN( u2_u6_u3_n165 ) );
  INV_X1 u2_u6_u3_U21 (.A( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n170 ) );
  NAND2_X1 u2_u6_u3_U22 (.A1( u2_u6_u3_n107 ) , .A2( u2_u6_u3_n108 ) , .ZN( u2_u6_u3_n140 ) );
  NAND2_X1 u2_u6_u3_U23 (.ZN( u2_u6_u3_n117 ) , .A1( u2_u6_u3_n124 ) , .A2( u2_u6_u3_n148 ) );
  NAND2_X1 u2_u6_u3_U24 (.ZN( u2_u6_u3_n143 ) , .A1( u2_u6_u3_n165 ) , .A2( u2_u6_u3_n167 ) );
  INV_X1 u2_u6_u3_U25 (.A( u2_u6_u3_n130 ) , .ZN( u2_u6_u3_n177 ) );
  INV_X1 u2_u6_u3_U26 (.A( u2_u6_u3_n128 ) , .ZN( u2_u6_u3_n176 ) );
  INV_X1 u2_u6_u3_U27 (.A( u2_u6_u3_n155 ) , .ZN( u2_u6_u3_n174 ) );
  AOI22_X1 u2_u6_u3_U28 (.B1( u2_u6_u3_n115 ) , .A2( u2_u6_u3_n116 ) , .ZN( u2_u6_u3_n123 ) , .B2( u2_u6_u3_n133 ) , .A1( u2_u6_u3_n169 ) );
  NAND2_X1 u2_u6_u3_U29 (.ZN( u2_u6_u3_n116 ) , .A2( u2_u6_u3_n151 ) , .A1( u2_u6_u3_n182 ) );
  INV_X1 u2_u6_u3_U3 (.A( u2_u6_u3_n129 ) , .ZN( u2_u6_u3_n183 ) );
  INV_X1 u2_u6_u3_U30 (.A( u2_u6_u3_n139 ) , .ZN( u2_u6_u3_n185 ) );
  NOR2_X1 u2_u6_u3_U31 (.ZN( u2_u6_u3_n135 ) , .A2( u2_u6_u3_n141 ) , .A1( u2_u6_u3_n169 ) );
  OAI222_X1 u2_u6_u3_U32 (.C2( u2_u6_u3_n107 ) , .A2( u2_u6_u3_n108 ) , .B1( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n138 ) , .B2( u2_u6_u3_n146 ) , .C1( u2_u6_u3_n154 ) , .A1( u2_u6_u3_n164 ) );
  NOR4_X1 u2_u6_u3_U33 (.A4( u2_u6_u3_n157 ) , .A3( u2_u6_u3_n158 ) , .A2( u2_u6_u3_n159 ) , .A1( u2_u6_u3_n160 ) , .ZN( u2_u6_u3_n161 ) );
  AOI21_X1 u2_u6_u3_U34 (.B2( u2_u6_u3_n152 ) , .B1( u2_u6_u3_n153 ) , .ZN( u2_u6_u3_n158 ) , .A( u2_u6_u3_n164 ) );
  AOI21_X1 u2_u6_u3_U35 (.A( u2_u6_u3_n154 ) , .B2( u2_u6_u3_n155 ) , .B1( u2_u6_u3_n156 ) , .ZN( u2_u6_u3_n157 ) );
  AOI21_X1 u2_u6_u3_U36 (.A( u2_u6_u3_n149 ) , .B2( u2_u6_u3_n150 ) , .B1( u2_u6_u3_n151 ) , .ZN( u2_u6_u3_n159 ) );
  AOI211_X1 u2_u6_u3_U37 (.ZN( u2_u6_u3_n109 ) , .A( u2_u6_u3_n119 ) , .C2( u2_u6_u3_n129 ) , .B( u2_u6_u3_n138 ) , .C1( u2_u6_u3_n141 ) );
  AOI211_X1 u2_u6_u3_U38 (.B( u2_u6_u3_n119 ) , .A( u2_u6_u3_n120 ) , .C2( u2_u6_u3_n121 ) , .ZN( u2_u6_u3_n122 ) , .C1( u2_u6_u3_n179 ) );
  INV_X1 u2_u6_u3_U39 (.A( u2_u6_u3_n156 ) , .ZN( u2_u6_u3_n179 ) );
  INV_X1 u2_u6_u3_U4 (.A( u2_u6_u3_n140 ) , .ZN( u2_u6_u3_n182 ) );
  OAI22_X1 u2_u6_u3_U40 (.B1( u2_u6_u3_n118 ) , .ZN( u2_u6_u3_n120 ) , .A1( u2_u6_u3_n135 ) , .B2( u2_u6_u3_n154 ) , .A2( u2_u6_u3_n178 ) );
  AND3_X1 u2_u6_u3_U41 (.ZN( u2_u6_u3_n118 ) , .A2( u2_u6_u3_n124 ) , .A1( u2_u6_u3_n144 ) , .A3( u2_u6_u3_n152 ) );
  INV_X1 u2_u6_u3_U42 (.A( u2_u6_u3_n121 ) , .ZN( u2_u6_u3_n164 ) );
  NAND2_X1 u2_u6_u3_U43 (.ZN( u2_u6_u3_n133 ) , .A1( u2_u6_u3_n154 ) , .A2( u2_u6_u3_n164 ) );
  OAI211_X1 u2_u6_u3_U44 (.B( u2_u6_u3_n127 ) , .ZN( u2_u6_u3_n139 ) , .C1( u2_u6_u3_n150 ) , .C2( u2_u6_u3_n154 ) , .A( u2_u6_u3_n184 ) );
  INV_X1 u2_u6_u3_U45 (.A( u2_u6_u3_n125 ) , .ZN( u2_u6_u3_n184 ) );
  AOI221_X1 u2_u6_u3_U46 (.A( u2_u6_u3_n126 ) , .ZN( u2_u6_u3_n127 ) , .C2( u2_u6_u3_n132 ) , .C1( u2_u6_u3_n169 ) , .B2( u2_u6_u3_n170 ) , .B1( u2_u6_u3_n174 ) );
  OAI22_X1 u2_u6_u3_U47 (.A1( u2_u6_u3_n124 ) , .ZN( u2_u6_u3_n125 ) , .B2( u2_u6_u3_n145 ) , .A2( u2_u6_u3_n165 ) , .B1( u2_u6_u3_n167 ) );
  NOR2_X1 u2_u6_u3_U48 (.A1( u2_u6_u3_n113 ) , .ZN( u2_u6_u3_n131 ) , .A2( u2_u6_u3_n154 ) );
  NAND2_X1 u2_u6_u3_U49 (.A1( u2_u6_u3_n103 ) , .ZN( u2_u6_u3_n150 ) , .A2( u2_u6_u3_n99 ) );
  INV_X1 u2_u6_u3_U5 (.A( u2_u6_u3_n117 ) , .ZN( u2_u6_u3_n178 ) );
  NAND2_X1 u2_u6_u3_U50 (.A2( u2_u6_u3_n102 ) , .ZN( u2_u6_u3_n155 ) , .A1( u2_u6_u3_n97 ) );
  INV_X1 u2_u6_u3_U51 (.A( u2_u6_u3_n141 ) , .ZN( u2_u6_u3_n167 ) );
  AOI21_X1 u2_u6_u3_U52 (.B2( u2_u6_u3_n114 ) , .B1( u2_u6_u3_n146 ) , .A( u2_u6_u3_n154 ) , .ZN( u2_u6_u3_n94 ) );
  AOI21_X1 u2_u6_u3_U53 (.ZN( u2_u6_u3_n110 ) , .B2( u2_u6_u3_n142 ) , .B1( u2_u6_u3_n186 ) , .A( u2_u6_u3_n95 ) );
  INV_X1 u2_u6_u3_U54 (.A( u2_u6_u3_n145 ) , .ZN( u2_u6_u3_n186 ) );
  AOI21_X1 u2_u6_u3_U55 (.B1( u2_u6_u3_n124 ) , .A( u2_u6_u3_n149 ) , .B2( u2_u6_u3_n155 ) , .ZN( u2_u6_u3_n95 ) );
  INV_X1 u2_u6_u3_U56 (.A( u2_u6_u3_n149 ) , .ZN( u2_u6_u3_n169 ) );
  NAND2_X1 u2_u6_u3_U57 (.ZN( u2_u6_u3_n124 ) , .A1( u2_u6_u3_n96 ) , .A2( u2_u6_u3_n97 ) );
  NAND2_X1 u2_u6_u3_U58 (.A2( u2_u6_u3_n100 ) , .ZN( u2_u6_u3_n146 ) , .A1( u2_u6_u3_n96 ) );
  NAND2_X1 u2_u6_u3_U59 (.A1( u2_u6_u3_n101 ) , .ZN( u2_u6_u3_n145 ) , .A2( u2_u6_u3_n99 ) );
  AOI221_X1 u2_u6_u3_U6 (.A( u2_u6_u3_n131 ) , .C2( u2_u6_u3_n132 ) , .C1( u2_u6_u3_n133 ) , .ZN( u2_u6_u3_n134 ) , .B1( u2_u6_u3_n143 ) , .B2( u2_u6_u3_n177 ) );
  NAND2_X1 u2_u6_u3_U60 (.A1( u2_u6_u3_n100 ) , .ZN( u2_u6_u3_n156 ) , .A2( u2_u6_u3_n99 ) );
  NAND2_X1 u2_u6_u3_U61 (.A2( u2_u6_u3_n101 ) , .A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n148 ) );
  NAND2_X1 u2_u6_u3_U62 (.A1( u2_u6_u3_n100 ) , .A2( u2_u6_u3_n102 ) , .ZN( u2_u6_u3_n128 ) );
  NAND2_X1 u2_u6_u3_U63 (.A2( u2_u6_u3_n101 ) , .A1( u2_u6_u3_n102 ) , .ZN( u2_u6_u3_n152 ) );
  NAND2_X1 u2_u6_u3_U64 (.A2( u2_u6_u3_n101 ) , .ZN( u2_u6_u3_n114 ) , .A1( u2_u6_u3_n96 ) );
  NAND2_X1 u2_u6_u3_U65 (.ZN( u2_u6_u3_n107 ) , .A1( u2_u6_u3_n97 ) , .A2( u2_u6_u3_n99 ) );
  NAND2_X1 u2_u6_u3_U66 (.A2( u2_u6_u3_n100 ) , .A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n113 ) );
  NAND2_X1 u2_u6_u3_U67 (.A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n153 ) , .A2( u2_u6_u3_n97 ) );
  NAND2_X1 u2_u6_u3_U68 (.A2( u2_u6_u3_n103 ) , .A1( u2_u6_u3_n104 ) , .ZN( u2_u6_u3_n130 ) );
  NAND2_X1 u2_u6_u3_U69 (.A2( u2_u6_u3_n103 ) , .ZN( u2_u6_u3_n144 ) , .A1( u2_u6_u3_n96 ) );
  OAI22_X1 u2_u6_u3_U7 (.B2( u2_u6_u3_n147 ) , .A2( u2_u6_u3_n148 ) , .ZN( u2_u6_u3_n160 ) , .B1( u2_u6_u3_n165 ) , .A1( u2_u6_u3_n168 ) );
  NAND2_X1 u2_u6_u3_U70 (.A1( u2_u6_u3_n102 ) , .A2( u2_u6_u3_n103 ) , .ZN( u2_u6_u3_n108 ) );
  NOR2_X1 u2_u6_u3_U71 (.A2( u2_u6_X_19 ) , .A1( u2_u6_X_20 ) , .ZN( u2_u6_u3_n99 ) );
  NOR2_X1 u2_u6_u3_U72 (.A2( u2_u6_X_21 ) , .A1( u2_u6_X_24 ) , .ZN( u2_u6_u3_n103 ) );
  NOR2_X1 u2_u6_u3_U73 (.A2( u2_u6_X_24 ) , .A1( u2_u6_u3_n171 ) , .ZN( u2_u6_u3_n97 ) );
  NOR2_X1 u2_u6_u3_U74 (.A2( u2_u6_X_23 ) , .ZN( u2_u6_u3_n141 ) , .A1( u2_u6_u3_n166 ) );
  NOR2_X1 u2_u6_u3_U75 (.A2( u2_u6_X_19 ) , .A1( u2_u6_u3_n172 ) , .ZN( u2_u6_u3_n96 ) );
  NAND2_X1 u2_u6_u3_U76 (.A1( u2_u6_X_22 ) , .A2( u2_u6_X_23 ) , .ZN( u2_u6_u3_n154 ) );
  NAND2_X1 u2_u6_u3_U77 (.A1( u2_u6_X_23 ) , .ZN( u2_u6_u3_n149 ) , .A2( u2_u6_u3_n166 ) );
  NOR2_X1 u2_u6_u3_U78 (.A2( u2_u6_X_22 ) , .A1( u2_u6_X_23 ) , .ZN( u2_u6_u3_n121 ) );
  AND2_X1 u2_u6_u3_U79 (.A1( u2_u6_X_24 ) , .ZN( u2_u6_u3_n101 ) , .A2( u2_u6_u3_n171 ) );
  AND3_X1 u2_u6_u3_U8 (.A3( u2_u6_u3_n144 ) , .A2( u2_u6_u3_n145 ) , .A1( u2_u6_u3_n146 ) , .ZN( u2_u6_u3_n147 ) );
  AND2_X1 u2_u6_u3_U80 (.A1( u2_u6_X_19 ) , .ZN( u2_u6_u3_n102 ) , .A2( u2_u6_u3_n172 ) );
  AND2_X1 u2_u6_u3_U81 (.A1( u2_u6_X_21 ) , .A2( u2_u6_X_24 ) , .ZN( u2_u6_u3_n100 ) );
  AND2_X1 u2_u6_u3_U82 (.A2( u2_u6_X_19 ) , .A1( u2_u6_X_20 ) , .ZN( u2_u6_u3_n104 ) );
  INV_X1 u2_u6_u3_U83 (.A( u2_u6_X_22 ) , .ZN( u2_u6_u3_n166 ) );
  INV_X1 u2_u6_u3_U84 (.A( u2_u6_X_21 ) , .ZN( u2_u6_u3_n171 ) );
  INV_X1 u2_u6_u3_U85 (.A( u2_u6_X_20 ) , .ZN( u2_u6_u3_n172 ) );
  NAND4_X1 u2_u6_u3_U86 (.ZN( u2_out6_26 ) , .A4( u2_u6_u3_n109 ) , .A3( u2_u6_u3_n110 ) , .A2( u2_u6_u3_n111 ) , .A1( u2_u6_u3_n173 ) );
  INV_X1 u2_u6_u3_U87 (.ZN( u2_u6_u3_n173 ) , .A( u2_u6_u3_n94 ) );
  OAI21_X1 u2_u6_u3_U88 (.ZN( u2_u6_u3_n111 ) , .B2( u2_u6_u3_n117 ) , .A( u2_u6_u3_n133 ) , .B1( u2_u6_u3_n176 ) );
  NAND4_X1 u2_u6_u3_U89 (.ZN( u2_out6_20 ) , .A4( u2_u6_u3_n122 ) , .A3( u2_u6_u3_n123 ) , .A1( u2_u6_u3_n175 ) , .A2( u2_u6_u3_n180 ) );
  INV_X1 u2_u6_u3_U9 (.A( u2_u6_u3_n143 ) , .ZN( u2_u6_u3_n168 ) );
  INV_X1 u2_u6_u3_U90 (.A( u2_u6_u3_n126 ) , .ZN( u2_u6_u3_n180 ) );
  INV_X1 u2_u6_u3_U91 (.A( u2_u6_u3_n112 ) , .ZN( u2_u6_u3_n175 ) );
  NAND4_X1 u2_u6_u3_U92 (.ZN( u2_out6_1 ) , .A4( u2_u6_u3_n161 ) , .A3( u2_u6_u3_n162 ) , .A2( u2_u6_u3_n163 ) , .A1( u2_u6_u3_n185 ) );
  NAND2_X1 u2_u6_u3_U93 (.ZN( u2_u6_u3_n163 ) , .A2( u2_u6_u3_n170 ) , .A1( u2_u6_u3_n176 ) );
  AOI22_X1 u2_u6_u3_U94 (.B2( u2_u6_u3_n140 ) , .B1( u2_u6_u3_n141 ) , .A2( u2_u6_u3_n142 ) , .ZN( u2_u6_u3_n162 ) , .A1( u2_u6_u3_n177 ) );
  OR4_X1 u2_u6_u3_U95 (.ZN( u2_out6_10 ) , .A4( u2_u6_u3_n136 ) , .A3( u2_u6_u3_n137 ) , .A1( u2_u6_u3_n138 ) , .A2( u2_u6_u3_n139 ) );
  OAI222_X1 u2_u6_u3_U96 (.C1( u2_u6_u3_n128 ) , .ZN( u2_u6_u3_n137 ) , .B1( u2_u6_u3_n148 ) , .A2( u2_u6_u3_n150 ) , .B2( u2_u6_u3_n154 ) , .C2( u2_u6_u3_n164 ) , .A1( u2_u6_u3_n167 ) );
  OAI221_X1 u2_u6_u3_U97 (.A( u2_u6_u3_n134 ) , .B2( u2_u6_u3_n135 ) , .ZN( u2_u6_u3_n136 ) , .C1( u2_u6_u3_n149 ) , .B1( u2_u6_u3_n151 ) , .C2( u2_u6_u3_n183 ) );
  NAND3_X1 u2_u6_u3_U98 (.A1( u2_u6_u3_n114 ) , .ZN( u2_u6_u3_n115 ) , .A2( u2_u6_u3_n145 ) , .A3( u2_u6_u3_n153 ) );
  NAND3_X1 u2_u6_u3_U99 (.ZN( u2_u6_u3_n129 ) , .A2( u2_u6_u3_n144 ) , .A1( u2_u6_u3_n153 ) , .A3( u2_u6_u3_n182 ) );
  OAI22_X1 u2_uk_U153 (.ZN( u2_K7_19 ) , .B2( u2_uk_n1465 ) , .A2( u2_uk_n1475 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U194 (.ZN( u2_K7_24 ) , .A( u2_uk_n1083 ) );
  AOI22_X1 u2_uk_U195 (.B2( u2_uk_K_r5_18 ) , .A2( u2_uk_K_r5_40 ) , .ZN( u2_uk_n1083 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n208 ) );
  OAI22_X1 u2_uk_U242 (.ZN( u2_K16_48 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1200 ) , .A2( u2_uk_n1208 ) , .A1( u2_uk_n213 ) );
  OAI21_X1 u2_uk_U598 (.ZN( u2_K7_22 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1081 ) , .B2( u2_uk_n1468 ) );
  OAI22_X1 u2_uk_U648 (.ZN( u2_K16_45 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1217 ) , .A2( u2_uk_n1220 ) , .A1( u2_uk_n238 ) );
  INV_X1 u2_uk_U661 (.ZN( u2_K16_43 ) , .A( u2_uk_n963 ) );
  AOI22_X1 u2_uk_U662 (.B2( u2_uk_K_r14_16 ) , .A2( u2_uk_K_r14_9 ) , .B1( u2_uk_n118 ) , .A1( u2_uk_n161 ) , .ZN( u2_uk_n963 ) );
  OAI21_X1 u2_uk_U782 (.ZN( u2_K7_21 ) , .A( u2_uk_n1080 ) , .B2( u2_uk_n1496 ) , .B1( u2_uk_n231 ) );
  NAND2_X1 u2_uk_U783 (.A1( u2_uk_K_r5_19 ) , .ZN( u2_uk_n1080 ) , .A2( u2_uk_n129 ) );
  INV_X1 u2_uk_U826 (.ZN( u2_K7_20 ) , .A( u2_uk_n1079 ) );
  OAI22_X1 u2_uk_U922 (.ZN( u2_K16_46 ) , .B2( u2_uk_n1189 ) , .A2( u2_uk_n1223 ) , .B1( u2_uk_n217 ) , .A1( u2_uk_n94 ) );
  OAI21_X1 u2_uk_U977 (.ZN( u2_K7_23 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1082 ) , .B2( u2_uk_n1453 ) );
endmodule

