module aes_aes_die_2 ( sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, 
       sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa12_0, sa12_1, 
       sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa31_0, sa31_1, sa31_2, 
       sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, w3_24, w3_25, w3_26, w3_27, 
       w3_28, w3_29, w3_30, w3_31, sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, 
        sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa11_sr_0, sa11_sr_1, 
        sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, 
        sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, u0_subword_0, u0_subword_1, u0_subword_2, u0_subword_3, 
        u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7 );
  input sa01_0, sa01_1, sa01_2, sa01_3, sa01_4, sa01_5, sa01_6, sa01_7, sa02_0, 
        sa02_1, sa02_2, sa02_3, sa02_4, sa02_5, sa02_6, sa02_7, sa12_0, sa12_1, 
        sa12_2, sa12_3, sa12_4, sa12_5, sa12_6, sa12_7, sa31_0, sa31_1, sa31_2, 
        sa31_3, sa31_4, sa31_5, sa31_6, sa31_7, w3_24, w3_25, w3_26, w3_27, 
        w3_28, w3_29, w3_30, w3_31;
  output sa01_sr_0, sa01_sr_1, sa01_sr_2, sa01_sr_3, sa01_sr_4, sa01_sr_5, sa01_sr_6, sa01_sr_7, sa02_sr_0, 
        sa02_sr_1, sa02_sr_2, sa02_sr_3, sa02_sr_4, sa02_sr_5, sa02_sr_6, sa02_sr_7, sa11_sr_0, sa11_sr_1, 
        sa11_sr_2, sa11_sr_3, sa11_sr_4, sa11_sr_5, sa11_sr_6, sa11_sr_7, sa32_sr_0, sa32_sr_1, sa32_sr_2, 
        sa32_sr_3, sa32_sr_4, sa32_sr_5, sa32_sr_6, sa32_sr_7, u0_subword_0, u0_subword_1, u0_subword_2, u0_subword_3, 
        u0_subword_4, u0_subword_5, u0_subword_6, u0_subword_7;
  wire u0_u3_n41, u0_u3_n438, u0_u3_n439, u0_u3_n440, u0_u3_n441, u0_u3_n442, u0_u3_n443, u0_u3_n444, u0_u3_n445, 
       u0_u3_n446, u0_u3_n447, u0_u3_n448, u0_u3_n449, u0_u3_n450, u0_u3_n451, u0_u3_n452, u0_u3_n453, u0_u3_n454, 
       u0_u3_n455, u0_u3_n456, u0_u3_n457, u0_u3_n458, u0_u3_n459, u0_u3_n460, u0_u3_n461, u0_u3_n462, u0_u3_n463, 
       u0_u3_n464, u0_u3_n465, u0_u3_n466, u0_u3_n467, u0_u3_n468, u0_u3_n469, u0_u3_n470, u0_u3_n471, u0_u3_n472, 
       u0_u3_n473, u0_u3_n474, u0_u3_n475, u0_u3_n476, u0_u3_n477, u0_u3_n478, u0_u3_n479, u0_u3_n480, u0_u3_n481, 
       u0_u3_n482, u0_u3_n483, u0_u3_n484, u0_u3_n485, u0_u3_n486, u0_u3_n487, u0_u3_n488, u0_u3_n489, u0_u3_n490, 
       u0_u3_n491, u0_u3_n492, u0_u3_n493, u0_u3_n494, u0_u3_n495, u0_u3_n496, u0_u3_n497, u0_u3_n498, u0_u3_n499, 
       u0_u3_n500, u0_u3_n501, u0_u3_n502, u0_u3_n503, u0_u3_n504, u0_u3_n505, u0_u3_n506, u0_u3_n507, u0_u3_n508, 
       u0_u3_n509, u0_u3_n510, u0_u3_n511, u0_u3_n512, u0_u3_n513, u0_u3_n514, u0_u3_n515, u0_u3_n516, u0_u3_n517, 
       u0_u3_n518, u0_u3_n519, u0_u3_n520, u0_u3_n521, u0_u3_n522, u0_u3_n523, u0_u3_n524, u0_u3_n525, u0_u3_n526, 
       u0_u3_n527, u0_u3_n528, u0_u3_n529, u0_u3_n530, u0_u3_n531, u0_u3_n532, u0_u3_n533, u0_u3_n534, u0_u3_n535, 
       u0_u3_n536, u0_u3_n537, u0_u3_n538, u0_u3_n539, u0_u3_n540, u0_u3_n541, u0_u3_n542, u0_u3_n543, u0_u3_n544, 
       u0_u3_n545, u0_u3_n546, u0_u3_n547, u0_u3_n548, u0_u3_n549, u0_u3_n550, u0_u3_n551, u0_u3_n552, u0_u3_n553, 
       u0_u3_n554, u0_u3_n555, u0_u3_n556, u0_u3_n557, u0_u3_n558, u0_u3_n559, u0_u3_n560, u0_u3_n561, u0_u3_n562, 
       u0_u3_n563, u0_u3_n564, u0_u3_n565, u0_u3_n566, u0_u3_n567, u0_u3_n568, u0_u3_n569, u0_u3_n570, u0_u3_n571, 
       u0_u3_n572, u0_u3_n573, u0_u3_n574, u0_u3_n575, u0_u3_n576, u0_u3_n577, u0_u3_n578, u0_u3_n579, u0_u3_n580, 
       u0_u3_n581, u0_u3_n582, u0_u3_n583, u0_u3_n584, u0_u3_n585, u0_u3_n586, u0_u3_n587, u0_u3_n588, u0_u3_n589, 
       u0_u3_n590, u0_u3_n591, u0_u3_n592, u0_u3_n593, u0_u3_n594, u0_u3_n595, u0_u3_n596, u0_u3_n597, u0_u3_n598, 
       u0_u3_n599, u0_u3_n600, u0_u3_n601, u0_u3_n602, u0_u3_n603, u0_u3_n604, u0_u3_n605, u0_u3_n606, u0_u3_n607, 
       u0_u3_n608, u0_u3_n609, u0_u3_n610, u0_u3_n611, u0_u3_n612, u0_u3_n613, u0_u3_n614, u0_u3_n615, u0_u3_n616, 
       u0_u3_n617, u0_u3_n618, u0_u3_n619, u0_u3_n620, u0_u3_n621, u0_u3_n622, u0_u3_n623, u0_u3_n624, u0_u3_n625, 
       u0_u3_n626, u0_u3_n627, u0_u3_n628, u0_u3_n629, u0_u3_n630, u0_u3_n631, u0_u3_n632, u0_u3_n633, u0_u3_n634, 
       u0_u3_n635, u0_u3_n636, u0_u3_n637, u0_u3_n638, u0_u3_n639, u0_u3_n640, u0_u3_n641, u0_u3_n642, u0_u3_n643, 
       u0_u3_n644, u0_u3_n645, u0_u3_n646, u0_u3_n647, u0_u3_n648, u0_u3_n649, u0_u3_n650, u0_u3_n651, u0_u3_n652, 
       u0_u3_n653, u0_u3_n654, u0_u3_n655, u0_u3_n656, u0_u3_n657, u0_u3_n658, u0_u3_n659, u0_u3_n660, u0_u3_n661, 
       u0_u3_n662, u0_u3_n663, u0_u3_n664, u0_u3_n665, u0_u3_n666, u0_u3_n667, u0_u3_n668, u0_u3_n669, u0_u3_n670, 
       u0_u3_n671, u0_u3_n672, u0_u3_n673, u0_u3_n674, u0_u3_n675, u0_u3_n676, u0_u3_n677, u0_u3_n678, u0_u3_n679, 
       u0_u3_n680, u0_u3_n681, u0_u3_n682, u0_u3_n683, u0_u3_n684, u0_u3_n685, u0_u3_n686, u0_u3_n687, u0_u3_n688, 
       u0_u3_n689, u0_u3_n690, u0_u3_n691, u0_u3_n692, u0_u3_n693, u0_u3_n694, u0_u3_n695, u0_u3_n696, u0_u3_n697, 
       u0_u3_n698, u0_u3_n699, u0_u3_n700, u0_u3_n701, u0_u3_n702, u0_u3_n703, u0_u3_n704, u0_u3_n705, u0_u3_n706, 
       u0_u3_n707, u0_u3_n708, u0_u3_n709, u0_u3_n710, u0_u3_n711, u0_u3_n712, u0_u3_n713, u0_u3_n714, u0_u3_n715, 
       u0_u3_n716, u0_u3_n717, u0_u3_n718, u0_u3_n719, u0_u3_n720, u0_u3_n721, u0_u3_n722, u0_u3_n723, u0_u3_n724, 
       u0_u3_n725, u0_u3_n726, u0_u3_n727, u0_u3_n728, u0_u3_n729, u0_u3_n730, u0_u3_n731, u0_u3_n732, u0_u3_n733, 
       u0_u3_n734, u0_u3_n735, u0_u3_n736, u0_u3_n737, u0_u3_n738, u0_u3_n739, u0_u3_n740, u0_u3_n741, u0_u3_n742, 
       u0_u3_n743, u0_u3_n744, u0_u3_n745, u0_u3_n746, u0_u3_n747, u0_u3_n748, u0_u3_n749, u0_u3_n750, u0_u3_n751, 
       u0_u3_n752, u0_u3_n753, u0_u3_n754, u0_u3_n755, u0_u3_n756, u0_u3_n757, u0_u3_n758, u0_u3_n759, u0_u3_n760, 
       u0_u3_n761, u0_u3_n762, u0_u3_n763, u0_u3_n764, u0_u3_n765, u0_u3_n766, u0_u3_n767, u0_u3_n768, u0_u3_n769, 
       u0_u3_n770, u0_u3_n771, u0_u3_n772, u0_u3_n773, u0_u3_n774, u0_u3_n775, u0_u3_n776, u0_u3_n777, u0_u3_n778, 
       u0_u3_n779, u0_u3_n780, u0_u3_n781, u0_u3_n782, u0_u3_n783, u0_u3_n784, u0_u3_n785, u0_u3_n786, u0_u3_n787, 
       u0_u3_n788, u0_u3_n789, u0_u3_n790, u0_u3_n791, u0_u3_n792, u0_u3_n793, u0_u3_n794, u0_u3_n795, u0_u3_n796, 
       u0_u3_n797, u0_u3_n798, u0_u3_n799, u0_u3_n800, u0_u3_n801, u0_u3_n802, u0_u3_n803, u0_u3_n804, u0_u3_n805, 
       u0_u3_n806, u0_u3_n807, u0_u3_n808, u0_u3_n809, u0_u3_n810, u0_u3_n811, u0_u3_n812, u0_u3_n813, u0_u3_n814, 
       u0_u3_n815, u0_u3_n816, u0_u3_n817, u0_u3_n818, u0_u3_n819, u0_u3_n820, u0_u3_n821, u0_u3_n822, u0_u3_n823, 
       u0_u3_n824, u0_u3_n825, u0_u3_n826, u0_u3_n827, u0_u3_n828, u0_u3_n829, u0_u3_n830, u0_u3_n831, u0_u3_n832, 
       u0_u3_n833, u0_u3_n834, u0_u3_n835, u0_u3_n836, u0_u3_n837, u0_u3_n838, u0_u3_n839, u0_u3_n840, u0_u3_n841, 
       u0_u3_n842, u0_u3_n843, u0_u3_n844, u0_u3_n845, u0_u3_n846, u0_u3_n847, u0_u3_n848, u0_u3_n849, u0_u3_n850, 
       u0_u3_n851, u0_u3_n852, u0_u3_n853, u0_u3_n854, u0_u3_n855, u0_u3_n856, u0_u3_n857, u0_u3_n858, u0_u3_n859, 
       u0_u3_n860, u0_u3_n861, u0_u3_n862, u0_u3_n863, u0_u3_n864, u0_u3_n865, u0_u3_n866, u0_u3_n867, u0_u3_n868, 
       u0_u3_n869, u0_u3_n870, u0_u3_n871, u0_u3_n872, u0_u3_n873, u0_u3_n874, u0_u3_n875, u0_u3_n876, u0_u3_n877, 
       u0_u3_n878, us01_n438, us01_n439, us01_n440, us01_n441, us01_n442, us01_n443, us01_n444, us01_n445, 
       us01_n446, us01_n447, us01_n448, us01_n449, us01_n450, us01_n451, us01_n452, us01_n453, us01_n454, 
       us01_n455, us01_n456, us01_n457, us01_n458, us01_n459, us01_n460, us01_n461, us01_n462, us01_n463, 
       us01_n464, us01_n465, us01_n466, us01_n467, us01_n468, us01_n469, us01_n470, us01_n471, us01_n472, 
       us01_n473, us01_n474, us01_n475, us01_n476, us01_n477, us01_n478, us01_n479, us01_n480, us01_n481, 
       us01_n482, us01_n483, us01_n484, us01_n485, us01_n486, us01_n487, us01_n488, us01_n489, us01_n490, 
       us01_n491, us01_n492, us01_n493, us01_n494, us01_n495, us01_n496, us01_n497, us01_n498, us01_n499, 
       us01_n500, us01_n501, us01_n502, us01_n503, us01_n504, us01_n505, us01_n506, us01_n507, us01_n508, 
       us01_n509, us01_n510, us01_n511, us01_n512, us01_n513, us01_n514, us01_n515, us01_n516, us01_n517, 
       us01_n518, us01_n519, us01_n520, us01_n521, us01_n522, us01_n523, us01_n524, us01_n525, us01_n526, 
       us01_n527, us01_n528, us01_n529, us01_n530, us01_n531, us01_n532, us01_n533, us01_n534, us01_n535, 
       us01_n536, us01_n537, us01_n538, us01_n539, us01_n540, us01_n541, us01_n542, us01_n543, us01_n544, 
       us01_n545, us01_n546, us01_n547, us01_n548, us01_n549, us01_n550, us01_n551, us01_n552, us01_n553, 
       us01_n554, us01_n555, us01_n556, us01_n557, us01_n558, us01_n559, us01_n560, us01_n561, us01_n562, 
       us01_n563, us01_n564, us01_n565, us01_n566, us01_n567, us01_n568, us01_n569, us01_n570, us01_n571, 
       us01_n572, us01_n573, us01_n574, us01_n575, us01_n576, us01_n577, us01_n578, us01_n579, us01_n580, 
       us01_n581, us01_n582, us01_n583, us01_n584, us01_n585, us01_n586, us01_n587, us01_n588, us01_n589, 
       us01_n590, us01_n591, us01_n592, us01_n593, us01_n594, us01_n595, us01_n596, us01_n597, us01_n598, 
       us01_n599, us01_n600, us01_n601, us01_n602, us01_n603, us01_n604, us01_n605, us01_n606, us01_n607, 
       us01_n608, us01_n609, us01_n610, us01_n611, us01_n612, us01_n613, us01_n614, us01_n615, us01_n616, 
       us01_n617, us01_n618, us01_n619, us01_n620, us01_n621, us01_n622, us01_n623, us01_n624, us01_n625, 
       us01_n626, us01_n627, us01_n628, us01_n629, us01_n630, us01_n631, us01_n632, us01_n633, us01_n634, 
       us01_n635, us01_n636, us01_n637, us01_n638, us01_n639, us01_n640, us01_n641, us01_n642, us01_n643, 
       us01_n644, us01_n645, us01_n646, us01_n647, us01_n648, us01_n649, us01_n650, us01_n651, us01_n652, 
       us01_n653, us01_n654, us01_n655, us01_n656, us01_n657, us01_n658, us01_n659, us01_n660, us01_n661, 
       us01_n662, us01_n663, us01_n664, us01_n665, us01_n666, us01_n667, us01_n668, us01_n669, us01_n670, 
       us01_n671, us01_n672, us01_n673, us01_n674, us01_n675, us01_n676, us01_n677, us01_n678, us01_n679, 
       us01_n680, us01_n681, us01_n682, us01_n683, us01_n684, us01_n685, us01_n686, us01_n687, us01_n688, 
       us01_n689, us01_n690, us01_n691, us01_n692, us01_n693, us01_n694, us01_n695, us01_n696, us01_n697, 
       us01_n698, us01_n699, us01_n700, us01_n701, us01_n702, us01_n703, us01_n704, us01_n705, us01_n706, 
       us01_n707, us01_n708, us01_n709, us01_n710, us01_n711, us01_n712, us01_n713, us01_n714, us01_n715, 
       us01_n716, us01_n717, us01_n718, us01_n719, us01_n720, us01_n721, us01_n722, us01_n723, us01_n724, 
       us01_n725, us01_n726, us01_n727, us01_n728, us01_n729, us01_n730, us01_n731, us01_n732, us01_n733, 
       us01_n734, us01_n735, us01_n736, us01_n737, us01_n738, us01_n739, us01_n740, us01_n741, us01_n742, 
       us01_n743, us01_n744, us01_n745, us01_n746, us01_n747, us01_n748, us01_n749, us01_n750, us01_n751, 
       us01_n752, us01_n753, us01_n754, us01_n755, us01_n756, us01_n757, us01_n758, us01_n759, us01_n760, 
       us01_n761, us01_n762, us01_n763, us01_n764, us01_n765, us01_n766, us01_n767, us01_n768, us01_n769, 
       us01_n770, us01_n771, us01_n772, us01_n773, us01_n774, us01_n775, us01_n776, us01_n777, us01_n778, 
       us01_n779, us01_n780, us01_n781, us01_n782, us01_n783, us01_n784, us01_n785, us01_n786, us01_n787, 
       us01_n788, us01_n789, us01_n790, us01_n791, us01_n792, us01_n793, us01_n794, us01_n795, us01_n796, 
       us01_n797, us01_n798, us01_n799, us01_n800, us01_n801, us01_n802, us01_n803, us01_n804, us01_n805, 
       us01_n806, us01_n807, us01_n808, us01_n809, us01_n810, us01_n811, us01_n812, us01_n813, us01_n814, 
       us01_n815, us01_n816, us01_n817, us01_n818, us01_n819, us01_n820, us01_n821, us01_n822, us01_n823, 
       us01_n824, us01_n825, us01_n826, us01_n827, us01_n828, us01_n829, us01_n830, us01_n831, us01_n832, 
       us01_n833, us01_n834, us01_n835, us01_n836, us01_n837, us01_n838, us01_n839, us01_n840, us01_n841, 
       us01_n842, us01_n843, us01_n844, us01_n845, us01_n846, us01_n847, us01_n848, us01_n849, us01_n850, 
       us01_n851, us01_n852, us01_n853, us01_n854, us01_n855, us01_n856, us01_n857, us01_n858, us01_n859, 
       us01_n860, us01_n861, us01_n862, us01_n863, us01_n864, us01_n865, us01_n866, us01_n867, us01_n868, 
       us01_n869, us01_n870, us01_n871, us01_n872, us01_n873, us01_n874, us02_n438, us02_n439, us02_n440, 
       us02_n441, us02_n442, us02_n443, us02_n444, us02_n445, us02_n446, us02_n447, us02_n448, us02_n449, 
       us02_n450, us02_n451, us02_n452, us02_n453, us02_n454, us02_n455, us02_n456, us02_n457, us02_n458, 
       us02_n459, us02_n460, us02_n461, us02_n462, us02_n463, us02_n464, us02_n465, us02_n466, us02_n467, 
       us02_n468, us02_n469, us02_n470, us02_n471, us02_n472, us02_n473, us02_n474, us02_n475, us02_n476, 
       us02_n477, us02_n478, us02_n479, us02_n480, us02_n481, us02_n482, us02_n483, us02_n484, us02_n485, 
       us02_n486, us02_n487, us02_n488, us02_n489, us02_n490, us02_n491, us02_n492, us02_n493, us02_n494, 
       us02_n495, us02_n496, us02_n497, us02_n498, us02_n499, us02_n500, us02_n501, us02_n502, us02_n503, 
       us02_n504, us02_n505, us02_n506, us02_n507, us02_n508, us02_n509, us02_n510, us02_n511, us02_n512, 
       us02_n513, us02_n514, us02_n515, us02_n516, us02_n517, us02_n518, us02_n519, us02_n520, us02_n521, 
       us02_n522, us02_n523, us02_n524, us02_n525, us02_n526, us02_n527, us02_n528, us02_n529, us02_n530, 
       us02_n531, us02_n532, us02_n533, us02_n534, us02_n535, us02_n536, us02_n537, us02_n538, us02_n539, 
       us02_n540, us02_n541, us02_n542, us02_n543, us02_n544, us02_n545, us02_n546, us02_n547, us02_n548, 
       us02_n549, us02_n550, us02_n551, us02_n552, us02_n553, us02_n554, us02_n555, us02_n556, us02_n557, 
       us02_n558, us02_n559, us02_n560, us02_n561, us02_n562, us02_n563, us02_n564, us02_n565, us02_n566, 
       us02_n567, us02_n568, us02_n569, us02_n570, us02_n571, us02_n572, us02_n573, us02_n574, us02_n575, 
       us02_n576, us02_n577, us02_n578, us02_n579, us02_n580, us02_n581, us02_n582, us02_n583, us02_n584, 
       us02_n585, us02_n586, us02_n587, us02_n588, us02_n589, us02_n590, us02_n591, us02_n592, us02_n593, 
       us02_n594, us02_n595, us02_n596, us02_n597, us02_n598, us02_n599, us02_n600, us02_n601, us02_n602, 
       us02_n603, us02_n604, us02_n605, us02_n606, us02_n607, us02_n608, us02_n609, us02_n610, us02_n611, 
       us02_n612, us02_n613, us02_n614, us02_n615, us02_n616, us02_n617, us02_n618, us02_n619, us02_n620, 
       us02_n621, us02_n622, us02_n623, us02_n624, us02_n625, us02_n626, us02_n627, us02_n628, us02_n629, 
       us02_n630, us02_n631, us02_n632, us02_n633, us02_n634, us02_n635, us02_n636, us02_n637, us02_n638, 
       us02_n639, us02_n640, us02_n641, us02_n642, us02_n643, us02_n644, us02_n645, us02_n646, us02_n647, 
       us02_n648, us02_n649, us02_n650, us02_n651, us02_n652, us02_n653, us02_n654, us02_n655, us02_n656, 
       us02_n657, us02_n658, us02_n659, us02_n660, us02_n661, us02_n662, us02_n663, us02_n664, us02_n665, 
       us02_n666, us02_n667, us02_n668, us02_n669, us02_n670, us02_n671, us02_n672, us02_n673, us02_n674, 
       us02_n675, us02_n676, us02_n677, us02_n678, us02_n679, us02_n680, us02_n681, us02_n682, us02_n683, 
       us02_n684, us02_n685, us02_n686, us02_n687, us02_n688, us02_n689, us02_n690, us02_n691, us02_n692, 
       us02_n693, us02_n694, us02_n695, us02_n696, us02_n697, us02_n698, us02_n699, us02_n700, us02_n701, 
       us02_n702, us02_n703, us02_n704, us02_n705, us02_n706, us02_n707, us02_n708, us02_n709, us02_n710, 
       us02_n711, us02_n712, us02_n713, us02_n714, us02_n715, us02_n716, us02_n717, us02_n718, us02_n719, 
       us02_n720, us02_n721, us02_n722, us02_n723, us02_n724, us02_n725, us02_n726, us02_n727, us02_n728, 
       us02_n729, us02_n730, us02_n731, us02_n732, us02_n733, us02_n734, us02_n735, us02_n736, us02_n737, 
       us02_n738, us02_n739, us02_n740, us02_n741, us02_n742, us02_n743, us02_n744, us02_n745, us02_n746, 
       us02_n747, us02_n748, us02_n749, us02_n750, us02_n751, us02_n752, us02_n753, us02_n754, us02_n755, 
       us02_n756, us02_n757, us02_n758, us02_n759, us02_n760, us02_n761, us02_n762, us02_n763, us02_n764, 
       us02_n765, us02_n766, us02_n767, us02_n768, us02_n769, us02_n770, us02_n771, us02_n772, us02_n773, 
       us02_n774, us02_n775, us02_n776, us02_n777, us02_n778, us02_n779, us02_n780, us02_n781, us02_n782, 
       us02_n783, us02_n784, us02_n785, us02_n786, us02_n787, us02_n788, us02_n789, us02_n790, us02_n791, 
       us02_n792, us02_n793, us02_n794, us02_n795, us02_n796, us02_n797, us02_n798, us02_n799, us02_n800, 
       us02_n801, us02_n802, us02_n803, us02_n804, us02_n805, us02_n806, us02_n807, us02_n808, us02_n809, 
       us02_n810, us02_n811, us02_n812, us02_n813, us02_n814, us02_n815, us02_n816, us02_n817, us02_n818, 
       us02_n819, us02_n820, us02_n821, us02_n822, us02_n823, us02_n824, us02_n825, us02_n826, us02_n827, 
       us02_n828, us02_n829, us02_n830, us02_n831, us02_n832, us02_n833, us02_n834, us02_n835, us02_n836, 
       us02_n837, us02_n838, us02_n839, us02_n840, us02_n841, us02_n842, us02_n843, us02_n844, us02_n845, 
       us02_n846, us02_n847, us02_n848, us02_n849, us02_n850, us02_n851, us02_n852, us02_n853, us02_n854, 
       us02_n855, us02_n856, us02_n857, us02_n858, us02_n859, us02_n860, us02_n861, us02_n862, us02_n863, 
       us02_n864, us02_n865, us02_n866, us02_n867, us02_n868, us02_n869, us02_n870, us02_n871, us02_n872, 
       us02_n873, us02_n874, us02_n875, us12_n438, us12_n439, us12_n440, us12_n441, us12_n442, us12_n443, 
       us12_n444, us12_n445, us12_n446, us12_n447, us12_n448, us12_n449, us12_n450, us12_n451, us12_n452, 
       us12_n453, us12_n454, us12_n455, us12_n456, us12_n457, us12_n458, us12_n459, us12_n460, us12_n461, 
       us12_n462, us12_n463, us12_n464, us12_n465, us12_n466, us12_n467, us12_n468, us12_n469, us12_n470, 
       us12_n471, us12_n472, us12_n473, us12_n474, us12_n475, us12_n476, us12_n477, us12_n478, us12_n479, 
       us12_n480, us12_n481, us12_n482, us12_n483, us12_n484, us12_n485, us12_n486, us12_n487, us12_n488, 
       us12_n489, us12_n490, us12_n491, us12_n492, us12_n493, us12_n494, us12_n495, us12_n496, us12_n497, 
       us12_n498, us12_n499, us12_n500, us12_n501, us12_n502, us12_n503, us12_n504, us12_n505, us12_n506, 
       us12_n507, us12_n508, us12_n509, us12_n510, us12_n511, us12_n512, us12_n513, us12_n514, us12_n515, 
       us12_n516, us12_n517, us12_n518, us12_n519, us12_n520, us12_n521, us12_n522, us12_n523, us12_n524, 
       us12_n525, us12_n526, us12_n527, us12_n528, us12_n529, us12_n530, us12_n531, us12_n532, us12_n533, 
       us12_n534, us12_n535, us12_n536, us12_n537, us12_n538, us12_n539, us12_n540, us12_n541, us12_n542, 
       us12_n543, us12_n544, us12_n545, us12_n546, us12_n547, us12_n548, us12_n549, us12_n550, us12_n551, 
       us12_n552, us12_n553, us12_n554, us12_n555, us12_n556, us12_n557, us12_n558, us12_n559, us12_n560, 
       us12_n561, us12_n562, us12_n563, us12_n564, us12_n565, us12_n566, us12_n567, us12_n568, us12_n569, 
       us12_n570, us12_n571, us12_n572, us12_n573, us12_n574, us12_n575, us12_n576, us12_n577, us12_n578, 
       us12_n579, us12_n580, us12_n581, us12_n582, us12_n583, us12_n584, us12_n585, us12_n586, us12_n587, 
       us12_n588, us12_n589, us12_n590, us12_n591, us12_n592, us12_n593, us12_n594, us12_n595, us12_n596, 
       us12_n597, us12_n598, us12_n599, us12_n600, us12_n601, us12_n602, us12_n603, us12_n604, us12_n605, 
       us12_n606, us12_n607, us12_n608, us12_n609, us12_n610, us12_n611, us12_n612, us12_n613, us12_n614, 
       us12_n615, us12_n616, us12_n617, us12_n618, us12_n619, us12_n620, us12_n621, us12_n622, us12_n623, 
       us12_n624, us12_n625, us12_n626, us12_n627, us12_n628, us12_n629, us12_n630, us12_n631, us12_n632, 
       us12_n633, us12_n634, us12_n635, us12_n636, us12_n637, us12_n638, us12_n639, us12_n640, us12_n641, 
       us12_n642, us12_n643, us12_n644, us12_n645, us12_n646, us12_n647, us12_n648, us12_n649, us12_n650, 
       us12_n651, us12_n652, us12_n653, us12_n654, us12_n655, us12_n656, us12_n657, us12_n658, us12_n659, 
       us12_n660, us12_n661, us12_n662, us12_n663, us12_n664, us12_n665, us12_n666, us12_n667, us12_n668, 
       us12_n669, us12_n670, us12_n671, us12_n672, us12_n673, us12_n674, us12_n675, us12_n676, us12_n677, 
       us12_n678, us12_n679, us12_n680, us12_n681, us12_n682, us12_n683, us12_n684, us12_n685, us12_n686, 
       us12_n687, us12_n688, us12_n689, us12_n690, us12_n691, us12_n692, us12_n693, us12_n694, us12_n695, 
       us12_n696, us12_n697, us12_n698, us12_n699, us12_n700, us12_n701, us12_n702, us12_n703, us12_n704, 
       us12_n705, us12_n706, us12_n707, us12_n708, us12_n709, us12_n710, us12_n711, us12_n712, us12_n713, 
       us12_n714, us12_n715, us12_n716, us12_n717, us12_n718, us12_n719, us12_n720, us12_n721, us12_n722, 
       us12_n723, us12_n724, us12_n725, us12_n726, us12_n727, us12_n728, us12_n729, us12_n730, us12_n731, 
       us12_n732, us12_n733, us12_n734, us12_n735, us12_n736, us12_n737, us12_n738, us12_n739, us12_n740, 
       us12_n741, us12_n742, us12_n743, us12_n744, us12_n745, us12_n746, us12_n747, us12_n748, us12_n749, 
       us12_n750, us12_n751, us12_n752, us12_n753, us12_n754, us12_n755, us12_n756, us12_n757, us12_n758, 
       us12_n759, us12_n760, us12_n761, us12_n762, us12_n763, us12_n764, us12_n765, us12_n766, us12_n767, 
       us12_n768, us12_n769, us12_n770, us12_n771, us12_n772, us12_n773, us12_n774, us12_n775, us12_n776, 
       us12_n777, us12_n778, us12_n779, us12_n780, us12_n781, us12_n782, us12_n783, us12_n784, us12_n785, 
       us12_n786, us12_n787, us12_n788, us12_n789, us12_n790, us12_n791, us12_n792, us12_n793, us12_n794, 
       us12_n795, us12_n796, us12_n797, us12_n798, us12_n799, us12_n800, us12_n801, us12_n802, us12_n803, 
       us12_n804, us12_n805, us12_n806, us12_n807, us12_n808, us12_n809, us12_n810, us12_n811, us12_n812, 
       us12_n813, us12_n814, us12_n815, us12_n816, us12_n817, us12_n818, us12_n819, us12_n820, us12_n821, 
       us12_n822, us12_n823, us12_n824, us12_n825, us12_n826, us12_n827, us12_n828, us12_n829, us12_n830, 
       us12_n831, us12_n832, us12_n833, us12_n834, us12_n835, us12_n836, us12_n837, us12_n838, us12_n839, 
       us12_n840, us12_n841, us12_n842, us12_n843, us12_n844, us12_n845, us12_n846, us12_n847, us12_n848, 
       us12_n849, us12_n850, us12_n851, us12_n852, us12_n853, us12_n854, us12_n855, us12_n856, us12_n857, 
       us12_n858, us12_n859, us12_n860, us12_n861, us12_n862, us12_n863, us12_n864, us12_n865, us12_n866, 
       us12_n867, us12_n868, us12_n869, us12_n870, us12_n871, us12_n872, us12_n873, us12_n874, us12_n875, 
       us12_n876, us31_n438, us31_n439, us31_n440, us31_n441, us31_n442, us31_n443, us31_n444, us31_n445, 
       us31_n446, us31_n447, us31_n448, us31_n449, us31_n450, us31_n451, us31_n452, us31_n453, us31_n454, 
       us31_n455, us31_n456, us31_n457, us31_n458, us31_n459, us31_n460, us31_n461, us31_n462, us31_n463, 
       us31_n464, us31_n465, us31_n466, us31_n467, us31_n468, us31_n469, us31_n470, us31_n471, us31_n472, 
       us31_n473, us31_n474, us31_n475, us31_n476, us31_n477, us31_n478, us31_n479, us31_n480, us31_n481, 
       us31_n482, us31_n483, us31_n484, us31_n485, us31_n486, us31_n487, us31_n488, us31_n489, us31_n490, 
       us31_n491, us31_n492, us31_n493, us31_n494, us31_n495, us31_n496, us31_n497, us31_n498, us31_n499, 
       us31_n500, us31_n501, us31_n502, us31_n503, us31_n504, us31_n505, us31_n506, us31_n507, us31_n508, 
       us31_n509, us31_n510, us31_n511, us31_n512, us31_n513, us31_n514, us31_n515, us31_n516, us31_n517, 
       us31_n518, us31_n519, us31_n520, us31_n521, us31_n522, us31_n523, us31_n524, us31_n525, us31_n526, 
       us31_n527, us31_n528, us31_n529, us31_n530, us31_n531, us31_n532, us31_n533, us31_n534, us31_n535, 
       us31_n536, us31_n537, us31_n538, us31_n539, us31_n540, us31_n541, us31_n542, us31_n543, us31_n544, 
       us31_n545, us31_n546, us31_n547, us31_n548, us31_n549, us31_n550, us31_n551, us31_n552, us31_n553, 
       us31_n554, us31_n555, us31_n556, us31_n557, us31_n558, us31_n559, us31_n560, us31_n561, us31_n562, 
       us31_n563, us31_n564, us31_n565, us31_n566, us31_n567, us31_n568, us31_n569, us31_n570, us31_n571, 
       us31_n572, us31_n573, us31_n574, us31_n575, us31_n576, us31_n577, us31_n578, us31_n579, us31_n580, 
       us31_n581, us31_n582, us31_n583, us31_n584, us31_n585, us31_n586, us31_n587, us31_n588, us31_n589, 
       us31_n590, us31_n591, us31_n592, us31_n593, us31_n594, us31_n595, us31_n596, us31_n597, us31_n598, 
       us31_n599, us31_n600, us31_n601, us31_n602, us31_n603, us31_n604, us31_n605, us31_n606, us31_n607, 
       us31_n608, us31_n609, us31_n610, us31_n611, us31_n612, us31_n613, us31_n614, us31_n615, us31_n616, 
       us31_n617, us31_n618, us31_n619, us31_n620, us31_n621, us31_n622, us31_n623, us31_n624, us31_n625, 
       us31_n626, us31_n627, us31_n628, us31_n629, us31_n630, us31_n631, us31_n632, us31_n633, us31_n634, 
       us31_n635, us31_n636, us31_n637, us31_n638, us31_n639, us31_n640, us31_n641, us31_n642, us31_n643, 
       us31_n644, us31_n645, us31_n646, us31_n647, us31_n648, us31_n649, us31_n650, us31_n651, us31_n652, 
       us31_n653, us31_n654, us31_n655, us31_n656, us31_n657, us31_n658, us31_n659, us31_n660, us31_n661, 
       us31_n662, us31_n663, us31_n664, us31_n665, us31_n666, us31_n667, us31_n668, us31_n669, us31_n670, 
       us31_n671, us31_n672, us31_n673, us31_n674, us31_n675, us31_n676, us31_n677, us31_n678, us31_n679, 
       us31_n680, us31_n681, us31_n682, us31_n683, us31_n684, us31_n685, us31_n686, us31_n687, us31_n688, 
       us31_n689, us31_n690, us31_n691, us31_n692, us31_n693, us31_n694, us31_n695, us31_n696, us31_n697, 
       us31_n698, us31_n699, us31_n700, us31_n701, us31_n702, us31_n703, us31_n704, us31_n705, us31_n706, 
       us31_n707, us31_n708, us31_n709, us31_n710, us31_n711, us31_n712, us31_n713, us31_n714, us31_n715, 
       us31_n716, us31_n717, us31_n718, us31_n719, us31_n720, us31_n721, us31_n722, us31_n723, us31_n724, 
       us31_n725, us31_n726, us31_n727, us31_n728, us31_n729, us31_n730, us31_n731, us31_n732, us31_n733, 
       us31_n734, us31_n735, us31_n736, us31_n737, us31_n738, us31_n739, us31_n740, us31_n741, us31_n742, 
       us31_n743, us31_n744, us31_n745, us31_n746, us31_n747, us31_n748, us31_n749, us31_n750, us31_n751, 
       us31_n752, us31_n753, us31_n754, us31_n755, us31_n756, us31_n757, us31_n758, us31_n759, us31_n760, 
       us31_n761, us31_n762, us31_n763, us31_n764, us31_n765, us31_n766, us31_n767, us31_n768, us31_n769, 
       us31_n770, us31_n771, us31_n772, us31_n773, us31_n774, us31_n775, us31_n776, us31_n777, us31_n778, 
       us31_n779, us31_n780, us31_n781, us31_n782, us31_n783, us31_n784, us31_n785, us31_n786, us31_n787, 
       us31_n788, us31_n789, us31_n790, us31_n791, us31_n792, us31_n793, us31_n794, us31_n795, us31_n796, 
       us31_n797, us31_n798, us31_n799, us31_n800, us31_n801, us31_n802, us31_n803, us31_n804, us31_n805, 
       us31_n806, us31_n807, us31_n808, us31_n809, us31_n810, us31_n811, us31_n812, us31_n813, us31_n814, 
       us31_n815, us31_n816, us31_n817, us31_n818, us31_n819, us31_n820, us31_n821, us31_n822, us31_n823, 
       us31_n824, us31_n825, us31_n826, us31_n827, us31_n828, us31_n829, us31_n830, us31_n831, us31_n832, 
       us31_n833, us31_n834, us31_n835, us31_n836, us31_n837, us31_n838, us31_n839, us31_n840, us31_n841, 
       us31_n842, us31_n843, us31_n844, us31_n845, us31_n846, us31_n847, us31_n848, us31_n849, us31_n850, 
       us31_n851, us31_n852, us31_n853, us31_n854, us31_n855, us31_n856, us31_n857, us31_n858, us31_n859, 
       us31_n860, us31_n861, us31_n862, us31_n863, us31_n864, us31_n865, us31_n866, us31_n867, us31_n868, 
       us31_n869, us31_n870, us31_n871, us31_n872, us31_n873, us31_n874, us31_n875,  us31_n876;
  NOR2_X1 u0_u3_U10 (.ZN( u0_u3_n578 ) , .A1( u0_u3_n625 ) , .A2( u0_u3_n748 ) );
  NOR2_X1 u0_u3_U100 (.ZN( u0_u3_n669 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U101 (.ZN( u0_u3_n535 ) , .A2( u0_u3_n752 ) , .A1( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U102 (.A2( u0_u3_n711 ) , .A1( u0_u3_n765 ) , .ZN( u0_u3_n797 ) );
  OAI22_X1 u0_u3_U103 (.B1( u0_u3_n493 ) , .ZN( u0_u3_n494 ) , .A1( u0_u3_n689 ) , .A2( u0_u3_n766 ) , .B2( u0_u3_n820 ) );
  NOR3_X1 u0_u3_U104 (.ZN( u0_u3_n493 ) , .A1( u0_u3_n785 ) , .A2( u0_u3_n852 ) , .A3( u0_u3_n865 ) );
  NOR2_X1 u0_u3_U105 (.ZN( u0_u3_n509 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n765 ) );
  NOR2_X1 u0_u3_U106 (.ZN( u0_u3_n520 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n806 ) );
  OAI21_X1 u0_u3_U107 (.ZN( u0_u3_n734 ) , .A( u0_u3_n836 ) , .B2( u0_u3_n854 ) , .B1( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U108 (.ZN( u0_u3_n604 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U109 (.A2( u0_u3_n711 ) , .A1( u0_u3_n753 ) , .ZN( u0_u3_n774 ) );
  NOR2_X1 u0_u3_U11 (.A1( u0_u3_n681 ) , .ZN( u0_u3_n696 ) , .A2( u0_u3_n810 ) );
  NOR2_X1 u0_u3_U110 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n670 ) , .A1( u0_u3_n753 ) );
  BUF_X2 u0_u3_U111 (.Z( u0_u3_n439 ) , .A( u0_u3_n794 ) );
  OAI21_X1 u0_u3_U112 (.ZN( u0_u3_n790 ) , .A( u0_u3_n841 ) , .B1( u0_u3_n865 ) , .B2( u0_u3_n875 ) );
  BUF_X2 u0_u3_U113 (.Z( u0_u3_n41 ) , .A( u0_u3_n700 ) );
  NOR2_X1 u0_u3_U114 (.ZN( u0_u3_n632 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U115 (.ZN( u0_u3_n512 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U116 (.ZN( u0_u3_n510 ) , .A1( u0_u3_n815 ) , .A2( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U117 (.ZN( u0_u3_n666 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U118 (.ZN( u0_u3_n546 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U119 (.ZN( u0_u3_n511 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n788 ) );
  INV_X1 u0_u3_U12 (.A( u0_u3_n683 ) , .ZN( u0_u3_n842 ) );
  NOR2_X1 u0_u3_U120 (.ZN( u0_u3_n547 ) , .A2( u0_u3_n788 ) , .A1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U121 (.ZN( u0_u3_n685 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U122 (.ZN( u0_u3_n572 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n765 ) , .A( u0_u3_n783 ) );
  NOR2_X1 u0_u3_U123 (.ZN( u0_u3_n714 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n766 ) );
  NOR2_X1 u0_u3_U124 (.ZN( u0_u3_n532 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n782 ) );
  AOI21_X1 u0_u3_U125 (.ZN( u0_u3_n518 ) , .A( u0_u3_n732 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U126 (.ZN( u0_u3_n617 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n815 ) );
  INV_X1 u0_u3_U127 (.A( u0_u3_n753 ) , .ZN( u0_u3_n844 ) );
  AOI21_X1 u0_u3_U128 (.ZN( u0_u3_n594 ) , .B2( u0_u3_n766 ) , .A( u0_u3_n788 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U129 (.ZN( u0_u3_n517 ) , .A( u0_u3_n782 ) , .B2( u0_u3_n795 ) , .B1( u0_u3_n815 ) );
  INV_X1 u0_u3_U13 (.A( u0_u3_n650 ) , .ZN( u0_u3_n872 ) );
  AOI21_X1 u0_u3_U130 (.B1( u0_u3_n689 ) , .ZN( u0_u3_n690 ) , .A( u0_u3_n731 ) , .B2( u0_u3_n764 ) );
  INV_X1 u0_u3_U131 (.A( u0_u3_n731 ) , .ZN( u0_u3_n854 ) );
  NOR2_X1 u0_u3_U132 (.ZN( u0_u3_n571 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n765 ) );
  INV_X1 u0_u3_U133 (.A( u0_u3_n795 ) , .ZN( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U134 (.A1( u0_u3_n752 ) , .ZN( u0_u3_n770 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U135 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n618 ) , .A1( u0_u3_n788 ) );
  AOI211_X1 u0_u3_U136 (.C2( u0_u3_n440 ) , .B( u0_u3_n626 ) , .A( u0_u3_n627 ) , .ZN( u0_u3_n638 ) , .C1( u0_u3_n865 ) );
  NOR4_X1 u0_u3_U137 (.A4( u0_u3_n632 ) , .A3( u0_u3_n633 ) , .A2( u0_u3_n634 ) , .A1( u0_u3_n635 ) , .ZN( u0_u3_n636 ) );
  NOR4_X1 u0_u3_U138 (.A4( u0_u3_n629 ) , .A3( u0_u3_n630 ) , .A2( u0_u3_n631 ) , .ZN( u0_u3_n637 ) , .A1( u0_u3_n667 ) );
  INV_X1 u0_u3_U139 (.A( u0_u3_n783 ) , .ZN( u0_u3_n852 ) );
  NOR4_X1 u0_u3_U14 (.A4( u0_u3_n547 ) , .A3( u0_u3_n548 ) , .A2( u0_u3_n549 ) , .A1( u0_u3_n550 ) , .ZN( u0_u3_n551 ) );
  OAI21_X1 u0_u3_U140 (.A( u0_u3_n701 ) , .ZN( u0_u3_n705 ) , .B2( u0_u3_n753 ) , .B1( u0_u3_n807 ) );
  OAI21_X1 u0_u3_U141 (.ZN( u0_u3_n701 ) , .B2( u0_u3_n836 ) , .B1( u0_u3_n840 ) , .A( u0_u3_n862 ) );
  INV_X1 u0_u3_U142 (.A( u0_u3_n732 ) , .ZN( u0_u3_n870 ) );
  NOR2_X1 u0_u3_U143 (.A2( u0_u3_n440 ) , .ZN( u0_u3_n628 ) , .A1( u0_u3_n841 ) );
  INV_X1 u0_u3_U144 (.A( u0_u3_n766 ) , .ZN( u0_u3_n868 ) );
  NOR2_X1 u0_u3_U145 (.ZN( u0_u3_n473 ) , .A2( u0_u3_n782 ) , .A1( u0_u3_n818 ) );
  INV_X1 u0_u3_U146 (.A( u0_u3_n440 ) , .ZN( u0_u3_n816 ) );
  INV_X1 u0_u3_U147 (.A( u0_u3_n820 ) , .ZN( u0_u3_n846 ) );
  NAND2_X1 u0_u3_U148 (.ZN( u0_u3_n717 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n783 ) );
  INV_X1 u0_u3_U149 (.A( u0_u3_n788 ) , .ZN( u0_u3_n848 ) );
  NOR4_X1 u0_u3_U15 (.A4( u0_u3_n448 ) , .A3( u0_u3_n449 ) , .A2( u0_u3_n519 ) , .A1( u0_u3_n544 ) , .ZN( u0_u3_n709 ) );
  AOI221_X1 u0_u3_U150 (.A( u0_u3_n767 ) , .ZN( u0_u3_n777 ) , .C2( u0_u3_n813 ) , .B2( u0_u3_n838 ) , .C1( u0_u3_n857 ) , .B1( u0_u3_n868 ) );
  INV_X1 u0_u3_U151 (.A( u0_u3_n764 ) , .ZN( u0_u3_n838 ) );
  AND2_X1 u0_u3_U152 (.ZN( u0_u3_n735 ) , .A1( u0_u3_n782 ) , .A2( u0_u3_n788 ) );
  AOI221_X1 u0_u3_U153 (.A( u0_u3_n453 ) , .ZN( u0_u3_n462 ) , .C2( u0_u3_n756 ) , .B1( u0_u3_n835 ) , .C1( u0_u3_n844 ) , .B2( u0_u3_n863 ) );
  AOI21_X1 u0_u3_U154 (.ZN( u0_u3_n453 ) , .B2( u0_u3_n795 ) , .A( u0_u3_n806 ) , .B1( u0_u3_n818 ) );
  AOI211_X1 u0_u3_U155 (.A( u0_u3_n591 ) , .ZN( u0_u3_n600 ) , .B( u0_u3_n624 ) , .C1( u0_u3_n847 ) , .C2( u0_u3_n857 ) );
  OAI221_X1 u0_u3_U156 (.A( u0_u3_n730 ) , .C2( u0_u3_n731 ) , .B2( u0_u3_n732 ) , .B1( u0_u3_n733 ) , .ZN( u0_u3_n740 ) , .C1( u0_u3_n820 ) );
  NAND2_X1 u0_u3_U157 (.A1( u0_u3_n444 ) , .A2( u0_u3_n467 ) , .ZN( u0_u3_n711 ) );
  NAND2_X1 u0_u3_U158 (.A2( u0_u3_n474 ) , .A1( u0_u3_n475 ) , .ZN( u0_u3_n820 ) );
  NAND2_X1 u0_u3_U159 (.A2( u0_u3_n463 ) , .A1( u0_u3_n468 ) , .ZN( u0_u3_n783 ) );
  OR3_X1 u0_u3_U16 (.ZN( u0_u3_n449 ) , .A1( u0_u3_n531 ) , .A3( u0_u3_n580 ) , .A2( u0_u3_n877 ) );
  NAND2_X1 u0_u3_U160 (.A1( u0_u3_n458 ) , .A2( u0_u3_n474 ) , .ZN( u0_u3_n806 ) );
  NAND2_X1 u0_u3_U161 (.A2( u0_u3_n451 ) , .A1( u0_u3_n463 ) , .ZN( u0_u3_n731 ) );
  NAND2_X1 u0_u3_U162 (.A1( u0_u3_n452 ) , .A2( u0_u3_n467 ) , .ZN( u0_u3_n727 ) );
  NAND2_X1 u0_u3_U163 (.A2( u0_u3_n457 ) , .A1( u0_u3_n475 ) , .ZN( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U164 (.ZN( u0_u3_n456 ) , .A1( u0_u3_n829 ) , .A2( u0_u3_n830 ) );
  NAND2_X1 u0_u3_U165 (.A2( u0_u3_n467 ) , .A1( u0_u3_n468 ) , .ZN( u0_u3_n815 ) );
  NAND2_X1 u0_u3_U166 (.A2( u0_u3_n451 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n732 ) );
  NAND2_X1 u0_u3_U167 (.A2( u0_u3_n452 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n766 ) );
  NAND2_X1 u0_u3_U168 (.A1( u0_u3_n454 ) , .A2( u0_u3_n474 ) , .ZN( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U169 (.A1( u0_u3_n456 ) , .A2( u0_u3_n464 ) , .ZN( u0_u3_n747 ) );
  OR4_X1 u0_u3_U17 (.A4( u0_u3_n445 ) , .A2( u0_u3_n446 ) , .A1( u0_u3_n447 ) , .ZN( u0_u3_n448 ) , .A3( u0_u3_n556 ) );
  NAND2_X1 u0_u3_U170 (.A2( u0_u3_n444 ) , .A1( u0_u3_n450 ) , .ZN( u0_u3_n787 ) );
  NAND2_X1 u0_u3_U171 (.A1( u0_u3_n454 ) , .A2( u0_u3_n457 ) , .ZN( u0_u3_n817 ) );
  NAND2_X1 u0_u3_U172 (.A1( u0_u3_n450 ) , .A2( u0_u3_n452 ) , .ZN( u0_u3_n808 ) );
  NAND2_X1 u0_u3_U173 (.A2( u0_u3_n456 ) , .A1( u0_u3_n458 ) , .ZN( u0_u3_n809 ) );
  NAND2_X1 u0_u3_U174 (.A1( u0_u3_n450 ) , .A2( u0_u3_n451 ) , .ZN( u0_u3_n789 ) );
  NAND2_X1 u0_u3_U175 (.A2( u0_u3_n464 ) , .A1( u0_u3_n465 ) , .ZN( u0_u3_n750 ) );
  NAND2_X1 u0_u3_U176 (.A1( u0_u3_n465 ) , .A2( u0_u3_n475 ) , .ZN( u0_u3_n791 ) );
  NAND2_X1 u0_u3_U177 (.A2( u0_u3_n457 ) , .A1( u0_u3_n458 ) , .ZN( u0_u3_n733 ) );
  NAND2_X1 u0_u3_U178 (.A1( u0_u3_n454 ) , .A2( u0_u3_n465 ) , .ZN( u0_u3_n793 ) );
  AND2_X1 u0_u3_U179 (.ZN( u0_u3_n440 ) , .A1( u0_u3_n457 ) , .A2( u0_u3_n464 ) );
  INV_X1 u0_u3_U18 (.A( u0_u3_n616 ) , .ZN( u0_u3_n877 ) );
  NOR2_X1 u0_u3_U180 (.ZN( u0_u3_n452 ) , .A1( u0_u3_n850 ) , .A2( w3_28 ) );
  NAND4_X1 u0_u3_U181 (.ZN( u0_subword_1 ) , .A4( u0_u3_n598 ) , .A3( u0_u3_n599 ) , .A2( u0_u3_n600 ) , .A1( u0_u3_n601 ) );
  AOI211_X1 u0_u3_U182 (.B( u0_u3_n592 ) , .A( u0_u3_n593 ) , .ZN( u0_u3_n599 ) , .C2( u0_u3_n814 ) , .C1( u0_u3_n836 ) );
  NOR4_X1 u0_u3_U183 (.A4( u0_u3_n594 ) , .A3( u0_u3_n595 ) , .A2( u0_u3_n596 ) , .A1( u0_u3_n597 ) , .ZN( u0_u3_n598 ) );
  NOR4_X1 u0_u3_U184 (.A4( u0_u3_n737 ) , .A3( u0_u3_n738 ) , .A2( u0_u3_n739 ) , .A1( u0_u3_n740 ) , .ZN( u0_u3_n741 ) );
  AOI211_X1 u0_u3_U185 (.B( u0_u3_n728 ) , .A( u0_u3_n729 ) , .ZN( u0_u3_n742 ) , .C1( u0_u3_n845 ) , .C2( u0_u3_n857 ) );
  AOI222_X1 u0_u3_U186 (.B2( u0_u3_n641 ) , .ZN( u0_u3_n647 ) , .B1( u0_u3_n843 ) , .A1( u0_u3_n844 ) , .C2( u0_u3_n848 ) , .C1( u0_u3_n865 ) , .A2( u0_u3_n867 ) );
  NOR4_X1 u0_u3_U187 (.A4( u0_u3_n642 ) , .A3( u0_u3_n643 ) , .A2( u0_u3_n644 ) , .A1( u0_u3_n645 ) , .ZN( u0_u3_n646 ) );
  AOI221_X1 u0_u3_U188 (.A( u0_u3_n784 ) , .ZN( u0_u3_n801 ) , .C2( u0_u3_n839 ) , .B2( u0_u3_n840 ) , .B1( u0_u3_n867 ) , .C1( u0_u3_n868 ) );
  NOR4_X1 u0_u3_U189 (.A4( u0_u3_n796 ) , .A3( u0_u3_n797 ) , .A2( u0_u3_n798 ) , .A1( u0_u3_n799 ) , .ZN( u0_u3_n800 ) );
  NOR4_X1 u0_u3_U19 (.ZN( u0_u3_n478 ) , .A1( u0_u3_n534 ) , .A3( u0_u3_n571 ) , .A4( u0_u3_n603 ) , .A2( u0_u3_n645 ) );
  NAND4_X1 u0_u3_U190 (.ZN( u0_subword_0 ) , .A4( u0_u3_n504 ) , .A3( u0_u3_n505 ) , .A2( u0_u3_n506 ) , .A1( u0_u3_n507 ) );
  NOR4_X1 u0_u3_U191 (.A4( u0_u3_n501 ) , .A3( u0_u3_n502 ) , .A2( u0_u3_n503 ) , .ZN( u0_u3_n504 ) , .A1( u0_u3_n530 ) );
  AOI221_X1 u0_u3_U192 (.A( u0_u3_n500 ) , .ZN( u0_u3_n505 ) , .B2( u0_u3_n845 ) , .C1( u0_u3_n848 ) , .C2( u0_u3_n862 ) , .B1( u0_u3_n864 ) );
  NOR4_X1 u0_u3_U193 (.A4( u0_u3_n703 ) , .A3( u0_u3_n704 ) , .A2( u0_u3_n705 ) , .A1( u0_u3_n706 ) , .ZN( u0_u3_n707 ) );
  NOR4_X1 u0_u3_U194 (.A3( u0_u3_n758 ) , .A2( u0_u3_n759 ) , .A1( u0_u3_n760 ) , .ZN( u0_u3_n761 ) , .A4( u0_u3_n871 ) );
  AOI211_X1 u0_u3_U195 (.B( u0_u3_n748 ) , .A( u0_u3_n749 ) , .ZN( u0_u3_n762 ) , .C1( u0_u3_n835 ) , .C2( u0_u3_n855 ) );
  NAND4_X1 u0_u3_U196 (.ZN( u0_subword_7 ) , .A4( u0_u3_n825 ) , .A3( u0_u3_n826 ) , .A2( u0_u3_n827 ) , .A1( u0_u3_n828 ) );
  NOR4_X1 u0_u3_U197 (.A4( u0_u3_n821 ) , .A3( u0_u3_n822 ) , .A2( u0_u3_n823 ) , .A1( u0_u3_n824 ) , .ZN( u0_u3_n825 ) );
  NAND2_X1 u0_u3_U198 (.A2( u0_u3_n464 ) , .A1( u0_u3_n474 ) , .ZN( u0_u3_n700 ) );
  NAND2_X1 u0_u3_U199 (.A2( u0_u3_n451 ) , .A1( u0_u3_n467 ) , .ZN( u0_u3_n818 ) );
  INV_X1 u0_u3_U20 (.A( u0_u3_n752 ) , .ZN( u0_u3_n865 ) );
  OAI21_X1 u0_u3_U200 (.B1( u0_u3_n756 ) , .ZN( u0_u3_n757 ) , .A( u0_u3_n847 ) , .B2( u0_u3_n870 ) );
  AOI221_X1 u0_u3_U201 (.A( u0_u3_n567 ) , .C2( u0_u3_n568 ) , .ZN( u0_u3_n577 ) , .B2( u0_u3_n847 ) , .B1( u0_u3_n854 ) , .C1( u0_u3_n855 ) );
  AOI222_X1 u0_u3_U202 (.ZN( u0_u3_n663 ) , .A2( u0_u3_n841 ) , .B1( u0_u3_n843 ) , .C2( u0_u3_n847 ) , .A1( u0_u3_n862 ) , .C1( u0_u3_n865 ) , .B2( u0_u3_n872 ) );
  AOI221_X1 u0_u3_U203 (.A( u0_u3_n713 ) , .ZN( u0_u3_n724 ) , .C2( u0_u3_n846 ) , .B2( u0_u3_n847 ) , .C1( u0_u3_n863 ) , .B1( u0_u3_n864 ) );
  NAND4_X1 u0_u3_U204 (.A4( u0_u3_n538 ) , .A3( u0_u3_n539 ) , .A2( u0_u3_n540 ) , .A1( u0_u3_n541 ) , .ZN( u0_u3_n625 ) );
  NOR4_X1 u0_u3_U205 (.A1( u0_u3_n534 ) , .ZN( u0_u3_n539 ) , .A2( u0_u3_n657 ) , .A4( u0_u3_n671 ) , .A3( u0_u3_n768 ) );
  NAND4_X1 u0_u3_U206 (.A4( u0_u3_n496 ) , .A3( u0_u3_n497 ) , .A1( u0_u3_n498 ) , .ZN( u0_u3_n805 ) , .A2( u0_u3_n869 ) );
  NOR4_X1 u0_u3_U207 (.A2( u0_u3_n494 ) , .A1( u0_u3_n495 ) , .ZN( u0_u3_n496 ) , .A3( u0_u3_n583 ) , .A4( u0_u3_n615 ) );
  NAND2_X1 u0_u3_U208 (.A1( u0_u3_n444 ) , .A2( u0_u3_n463 ) , .ZN( u0_u3_n702 ) );
  NAND2_X1 u0_u3_U209 (.A1( u0_u3_n455 ) , .A2( u0_u3_n468 ) , .ZN( u0_u3_n672 ) );
  AOI222_X1 u0_u3_U21 (.ZN( u0_u3_n566 ) , .B1( u0_u3_n833 ) , .C1( u0_u3_n843 ) , .A2( u0_u3_n845 ) , .A1( u0_u3_n856 ) , .B2( u0_u3_n865 ) , .C2( u0_u3_n875 ) );
  NAND4_X1 u0_u3_U210 (.A4( u0_u3_n563 ) , .A3( u0_u3_n564 ) , .A2( u0_u3_n565 ) , .A1( u0_u3_n566 ) , .ZN( u0_u3_n610 ) );
  NOR4_X1 u0_u3_U211 (.ZN( u0_u3_n564 ) , .A1( u0_u3_n656 ) , .A3( u0_u3_n664 ) , .A4( u0_u3_n688 ) , .A2( u0_u3_n771 ) );
  NOR2_X1 u0_u3_U212 (.ZN( u0_u3_n454 ) , .A1( u0_u3_n831 ) , .A2( u0_u3_n832 ) );
  INV_X1 u0_u3_U213 (.ZN( u0_u3_n831 ) , .A( w3_26 ) );
  NOR2_X1 u0_u3_U214 (.ZN( u0_u3_n710 ) , .A2( u0_u3_n779 ) , .A1( u0_u3_n803 ) );
  OAI21_X1 u0_u3_U215 (.A( u0_u3_n734 ) , .B1( u0_u3_n735 ) , .ZN( u0_u3_n739 ) , .B2( u0_u3_n808 ) );
  AOI21_X1 u0_u3_U216 (.ZN( u0_u3_n653 ) , .A( u0_u3_n782 ) , .B1( u0_u3_n795 ) , .B2( u0_u3_n808 ) );
  INV_X1 u0_u3_U217 (.A( u0_u3_n808 ) , .ZN( u0_u3_n862 ) );
  NOR2_X1 u0_u3_U218 (.ZN( u0_u3_n738 ) , .A2( u0_u3_n806 ) , .A1( u0_u3_n808 ) );
  NAND2_X1 u0_u3_U219 (.ZN( u0_u3_n756 ) , .A1( u0_u3_n766 ) , .A2( u0_u3_n808 ) );
  NOR4_X1 u0_u3_U22 (.ZN( u0_u3_n482 ) , .A1( u0_u3_n523 ) , .A4( u0_u3_n560 ) , .A3( u0_u3_n585 ) , .A2( u0_u3_n633 ) );
  NOR2_X1 u0_u3_U220 (.ZN( u0_u3_n559 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n808 ) );
  OAI221_X1 u0_u3_U221 (.A( u0_u3_n699 ) , .ZN( u0_u3_n706 ) , .C2( u0_u3_n787 ) , .C1( u0_u3_n788 ) , .B1( u0_u3_n789 ) , .B2( u0_u3_n809 ) );
  OAI222_X1 u0_u3_U222 (.B1( u0_u3_n41 ) , .ZN( u0_u3_n620 ) , .C1( u0_u3_n727 ) , .C2( u0_u3_n750 ) , .B2( u0_u3_n789 ) , .A2( u0_u3_n795 ) , .A1( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U223 (.A2( u0_u3_n444 ) , .A1( u0_u3_n455 ) , .ZN( u0_u3_n794 ) );
  OAI222_X1 u0_u3_U224 (.B2( u0_u3_n711 ) , .ZN( u0_u3_n712 ) , .C2( u0_u3_n727 ) , .B1( u0_u3_n750 ) , .A1( u0_u3_n809 ) , .C1( u0_u3_n817 ) , .A2( u0_u3_n818 ) );
  INV_X1 u0_u3_U225 (.A( u0_u3_n675 ) , .ZN( u0_u3_n861 ) );
  NOR2_X1 u0_u3_U226 (.ZN( u0_u3_n531 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U227 (.ZN( u0_u3_n529 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n753 ) );
  INV_X1 u0_u3_U228 (.A( u0_u3_n727 ) , .ZN( u0_u3_n858 ) );
  NOR2_X1 u0_u3_U229 (.ZN( u0_u3_n450 ) , .A2( u0_u3_n851 ) , .A1( u0_u3_n860 ) );
  NOR4_X1 u0_u3_U23 (.A4( u0_u3_n559 ) , .A3( u0_u3_n560 ) , .A2( u0_u3_n561 ) , .A1( u0_u3_n562 ) , .ZN( u0_u3_n563 ) );
  AOI222_X1 u0_u3_U230 (.ZN( u0_u3_n528 ) , .A1( u0_u3_n837 ) , .B2( u0_u3_n839 ) , .C1( u0_u3_n846 ) , .C2( u0_u3_n852 ) , .A2( u0_u3_n854 ) , .B1( u0_u3_n868 ) );
  NOR3_X1 u0_u3_U231 (.A2( u0_u3_n440 ) , .ZN( u0_u3_n443 ) , .A3( u0_u3_n839 ) , .A1( u0_u3_n848 ) );
  NAND2_X1 u0_u3_U232 (.ZN( u0_u3_n616 ) , .A2( u0_u3_n839 ) , .A1( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U233 (.ZN( u0_u3_n498 ) , .A1( u0_u3_n681 ) , .A2( u0_u3_n697 ) );
  AOI211_X1 u0_u3_U234 (.B( u0_u3_n697 ) , .A( u0_u3_n698 ) , .ZN( u0_u3_n708 ) , .C2( u0_u3_n834 ) , .C1( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U235 (.ZN( u0_u3_n586 ) , .A1( u0_u3_n795 ) , .A2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U236 (.ZN( u0_u3_n543 ) , .A( u0_u3_n766 ) , .B2( u0_u3_n782 ) , .B1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U237 (.ZN( u0_u3_n612 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U238 (.ZN( u0_u3_n718 ) , .A1( u0_u3_n808 ) , .A2( u0_u3_n820 ) );
  OAI21_X1 u0_u3_U239 (.A( u0_u3_n790 ) , .B2( u0_u3_n791 ) , .B1( u0_u3_n792 ) , .ZN( u0_u3_n798 ) );
  NOR4_X1 u0_u3_U24 (.A4( u0_u3_n555 ) , .A3( u0_u3_n556 ) , .A2( u0_u3_n557 ) , .A1( u0_u3_n558 ) , .ZN( u0_u3_n565 ) );
  AOI21_X1 u0_u3_U240 (.ZN( u0_u3_n642 ) , .B2( u0_u3_n752 ) , .A( u0_u3_n791 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U241 (.A( u0_u3_n736 ) , .ZN( u0_u3_n737 ) , .B2( u0_u3_n783 ) , .B1( u0_u3_n795 ) );
  AOI21_X1 u0_u3_U242 (.B2( u0_u3_n766 ) , .ZN( u0_u3_n767 ) , .A( u0_u3_n791 ) , .B1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U243 (.ZN( u0_u3_n521 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U244 (.ZN( u0_u3_n487 ) , .A1( u0_u3_n791 ) , .A2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U245 (.ZN( u0_u3_n537 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n791 ) );
  INV_X1 u0_u3_U246 (.A( u0_u3_n791 ) , .ZN( u0_u3_n847 ) );
  OAI22_X1 u0_u3_U247 (.B2( u0_u3_n782 ) , .B1( u0_u3_n783 ) , .ZN( u0_u3_n784 ) , .A2( u0_u3_n817 ) , .A1( u0_u3_n818 ) );
  AOI21_X1 u0_u3_U248 (.ZN( u0_u3_n501 ) , .A( u0_u3_n727 ) , .B2( u0_u3_n765 ) , .B1( u0_u3_n817 ) );
  NAND4_X1 u0_u3_U249 (.A4( u0_u3_n482 ) , .A3( u0_u3_n483 ) , .A2( u0_u3_n484 ) , .A1( u0_u3_n485 ) , .ZN( u0_u3_n697 ) );
  NOR4_X1 u0_u3_U25 (.A4( u0_u3_n771 ) , .A3( u0_u3_n772 ) , .A2( u0_u3_n773 ) , .A1( u0_u3_n774 ) , .ZN( u0_u3_n775 ) );
  AOI21_X1 u0_u3_U250 (.ZN( u0_u3_n542 ) , .B2( u0_u3_n815 ) , .A( u0_u3_n817 ) , .B1( u0_u3_n818 ) );
  NOR2_X1 u0_u3_U251 (.ZN( u0_u3_n523 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U252 (.ZN( u0_u3_n549 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n817 ) );
  INV_X1 u0_u3_U253 (.A( u0_u3_n817 ) , .ZN( u0_u3_n836 ) );
  NOR2_X1 u0_u3_U254 (.ZN( u0_u3_n548 ) , .A1( u0_u3_n752 ) , .A2( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U255 (.ZN( u0_u3_n560 ) , .A1( u0_u3_n795 ) , .A2( u0_u3_n817 ) );
  AOI21_X1 u0_u3_U256 (.A( u0_u3_n673 ) , .B1( u0_u3_n674 ) , .ZN( u0_u3_n675 ) , .B2( u0_u3_n858 ) );
  AOI22_X1 u0_u3_U257 (.A2( u0_u3_n785 ) , .ZN( u0_u3_n786 ) , .B2( u0_u3_n834 ) , .A1( u0_u3_n837 ) , .B1( u0_u3_n865 ) );
  AOI21_X1 u0_u3_U258 (.ZN( u0_u3_n643 ) , .B2( u0_u3_n750 ) , .A( u0_u3_n795 ) , .B1( u0_u3_n806 ) );
  NAND4_X1 u0_u3_U259 (.A4( u0_u3_n775 ) , .A3( u0_u3_n776 ) , .A2( u0_u3_n777 ) , .A1( u0_u3_n778 ) , .ZN( u0_u3_n804 ) );
  NOR3_X1 u0_u3_U26 (.A3( u0_u3_n768 ) , .A2( u0_u3_n769 ) , .A1( u0_u3_n770 ) , .ZN( u0_u3_n776 ) );
  OAI21_X1 u0_u3_U260 (.ZN( u0_u3_n466 ) , .B1( u0_u3_n812 ) , .A( u0_u3_n837 ) , .B2( u0_u3_n853 ) );
  NOR2_X1 u0_u3_U261 (.ZN( u0_u3_n659 ) , .A1( u0_u3_n750 ) , .A2( u0_u3_n783 ) );
  NOR2_X1 u0_u3_U262 (.ZN( u0_u3_n683 ) , .A2( u0_u3_n837 ) , .A1( u0_u3_n841 ) );
  NOR2_X1 u0_u3_U263 (.ZN( u0_u3_n764 ) , .A1( u0_u3_n836 ) , .A2( u0_u3_n837 ) );
  NOR2_X1 u0_u3_U264 (.ZN( u0_u3_n570 ) , .A1( u0_u3_n750 ) , .A2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U265 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n633 ) , .A1( u0_u3_n750 ) );
  INV_X1 u0_u3_U266 (.A( u0_u3_n750 ) , .ZN( u0_u3_n837 ) );
  NOR4_X1 u0_u3_U267 (.ZN( u0_u3_n488 ) , .A2( u0_u3_n536 ) , .A1( u0_u3_n561 ) , .A3( u0_u3_n634 ) , .A4( u0_u3_n721 ) );
  NAND4_X1 u0_u3_U268 (.A4( u0_u3_n488 ) , .A3( u0_u3_n489 ) , .A2( u0_u3_n490 ) , .A1( u0_u3_n491 ) , .ZN( u0_u3_n781 ) );
  AOI21_X1 u0_u3_U269 (.B1( u0_u3_n438 ) , .ZN( u0_u3_n592 ) , .B2( u0_u3_n702 ) , .A( u0_u3_n820 ) );
  NAND4_X1 u0_u3_U27 (.A4( u0_u3_n606 ) , .A3( u0_u3_n607 ) , .A2( u0_u3_n608 ) , .A1( u0_u3_n609 ) , .ZN( u0_u3_n725 ) );
  AOI21_X1 u0_u3_U270 (.B1( u0_u3_n702 ) , .ZN( u0_u3_n703 ) , .A( u0_u3_n735 ) , .B2( u0_u3_n766 ) );
  INV_X1 u0_u3_U271 (.A( u0_u3_n702 ) , .ZN( u0_u3_n855 ) );
  AOI21_X1 u0_u3_U272 (.ZN( u0_u3_n445 ) , .A( u0_u3_n702 ) , .B1( u0_u3_n736 ) , .B2( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U273 (.ZN( u0_u3_n686 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U274 (.ZN( u0_u3_n580 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n817 ) );
  NAND2_X1 u0_u3_U275 (.A1( u0_u3_n702 ) , .A2( u0_u3_n732 ) , .ZN( u0_u3_n785 ) );
  NOR3_X1 u0_u3_U276 (.A3( u0_u3_n744 ) , .A2( u0_u3_n745 ) , .A1( u0_u3_n746 ) , .ZN( u0_u3_n763 ) );
  OAI22_X1 u0_u3_U277 (.ZN( u0_u3_n492 ) , .A1( u0_u3_n727 ) , .B2( u0_u3_n731 ) , .B1( u0_u3_n733 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U278 (.ZN( u0_u3_n582 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n733 ) );
  NOR2_X1 u0_u3_U279 (.ZN( u0_u3_n536 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n733 ) );
  NOR3_X1 u0_u3_U28 (.A1( u0_u3_n602 ) , .ZN( u0_u3_n607 ) , .A3( u0_u3_n666 ) , .A2( u0_u3_n773 ) );
  AOI222_X1 u0_u3_U280 (.ZN( u0_u3_n608 ) , .B2( u0_u3_n674 ) , .B1( u0_u3_n756 ) , .C2( u0_u3_n834 ) , .A1( u0_u3_n836 ) , .A2( u0_u3_n864 ) , .C1( u0_u3_n865 ) );
  AOI221_X1 u0_u3_U281 (.A( u0_u3_n486 ) , .ZN( u0_u3_n491 ) , .B1( u0_u3_n834 ) , .C2( u0_u3_n846 ) , .C1( u0_u3_n854 ) , .B2( u0_u3_n864 ) );
  NOR2_X1 u0_u3_U282 (.ZN( u0_u3_n792 ) , .A2( u0_u3_n864 ) , .A1( u0_u3_n870 ) );
  NOR2_X1 u0_u3_U283 (.ZN( u0_u3_n464 ) , .A1( u0_u3_n832 ) , .A2( w3_26 ) );
  NOR2_X1 u0_u3_U284 (.ZN( u0_u3_n474 ) , .A1( u0_u3_n829 ) , .A2( w3_25 ) );
  AOI21_X1 u0_u3_U285 (.A( u0_u3_n439 ) , .ZN( u0_u3_n644 ) , .B1( u0_u3_n683 ) , .B2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U286 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n500 ) , .A( u0_u3_n782 ) , .B1( u0_u3_n807 ) );
  OAI22_X1 u0_u3_U287 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n698 ) , .A2( u0_u3_n733 ) , .A1( u0_u3_n783 ) , .B2( u0_u3_n820 ) );
  AOI21_X1 u0_u3_U288 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n567 ) , .B1( u0_u3_n727 ) , .A( u0_u3_n782 ) );
  AOI21_X1 u0_u3_U289 (.B2( u0_u3_n439 ) , .ZN( u0_u3_n446 ) , .B1( u0_u3_n792 ) , .A( u0_u3_n817 ) );
  NOR4_X1 u0_u3_U29 (.A3( u0_u3_n603 ) , .A2( u0_u3_n604 ) , .A1( u0_u3_n605 ) , .ZN( u0_u3_n606 ) , .A4( u0_u3_n658 ) );
  NOR2_X1 u0_u3_U290 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n667 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U291 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n558 ) , .A1( u0_u3_n753 ) );
  NOR2_X1 u0_u3_U292 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n562 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U293 (.A1( u0_u3_n439 ) , .ZN( u0_u3_n645 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U294 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n545 ) , .A1( u0_u3_n765 ) );
  INV_X1 u0_u3_U295 (.A( u0_u3_n794 ) , .ZN( u0_u3_n875 ) );
  NOR2_X1 u0_u3_U296 (.ZN( u0_u3_n463 ) , .A1( u0_u3_n851 ) , .A2( w3_31 ) );
  AOI21_X1 u0_u3_U297 (.B2( u0_u3_n439 ) , .A( u0_u3_n793 ) , .B1( u0_u3_n795 ) , .ZN( u0_u3_n796 ) );
  AOI222_X1 u0_u3_U298 (.C2( u0_u3_n812 ) , .B2( u0_u3_n813 ) , .A2( u0_u3_n814 ) , .ZN( u0_u3_n826 ) , .C1( u0_u3_n835 ) , .A1( u0_u3_n841 ) , .B1( u0_u3_n855 ) );
  AOI22_X1 u0_u3_U299 (.ZN( u0_u3_n730 ) , .B1( u0_u3_n835 ) , .A2( u0_u3_n840 ) , .A1( u0_u3_n865 ) , .B2( u0_u3_n868 ) );
  BUF_X1 u0_u3_U3 (.Z( u0_u3_n438 ) , .A( u0_u3_n818 ) );
  NOR4_X1 u0_u3_U30 (.A4( u0_u3_n487 ) , .ZN( u0_u3_n490 ) , .A1( u0_u3_n569 ) , .A2( u0_u3_n584 ) , .A3( u0_u3_n605 ) );
  AOI222_X1 u0_u3_U300 (.ZN( u0_u3_n516 ) , .C1( u0_u3_n835 ) , .B2( u0_u3_n839 ) , .A2( u0_u3_n845 ) , .C2( u0_u3_n864 ) , .B1( u0_u3_n865 ) , .A1( u0_u3_n868 ) );
  AOI222_X1 u0_u3_U301 (.ZN( u0_u3_n472 ) , .B1( u0_u3_n835 ) , .A1( u0_u3_n841 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n853 ) , .A2( u0_u3_n857 ) , .B2( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U302 (.A2( u0_u3_n438 ) , .ZN( u0_u3_n658 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U303 (.ZN( u0_u3_n715 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U304 (.ZN( u0_u3_n689 ) , .A1( u0_u3_n834 ) , .A2( u0_u3_n835 ) );
  NOR2_X1 u0_u3_U305 (.ZN( u0_u3_n524 ) , .A1( u0_u3_n793 ) , .A2( u0_u3_n815 ) );
  NOR2_X1 u0_u3_U306 (.ZN( u0_u3_n664 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U307 (.ZN( u0_u3_n736 ) , .A2( u0_u3_n835 ) , .A1( u0_u3_n847 ) );
  NOR2_X1 u0_u3_U308 (.ZN( u0_u3_n671 ) , .A2( u0_u3_n711 ) , .A1( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U309 (.ZN( u0_u3_n673 ) , .A1( u0_u3_n793 ) , .A2( u0_u3_n808 ) );
  NOR4_X1 u0_u3_U31 (.ZN( u0_u3_n489 ) , .A1( u0_u3_n510 ) , .A2( u0_u3_n522 ) , .A4( u0_u3_n549 ) , .A3( u0_u3_n614 ) );
  INV_X1 u0_u3_U310 (.A( u0_u3_n793 ) , .ZN( u0_u3_n835 ) );
  AOI21_X1 u0_u3_U311 (.B1( u0_u3_n438 ) , .ZN( u0_u3_n513 ) , .B2( u0_u3_n672 ) , .A( u0_u3_n733 ) );
  AOI21_X1 u0_u3_U312 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n629 ) , .B2( u0_u3_n672 ) , .A( u0_u3_n793 ) );
  INV_X1 u0_u3_U313 (.A( u0_u3_n672 ) , .ZN( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U314 (.ZN( u0_u3_n655 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n817 ) );
  NOR2_X1 u0_u3_U315 (.ZN( u0_u3_n631 ) , .A2( u0_u3_n672 ) , .A1( u0_u3_n788 ) );
  NOR2_X1 u0_u3_U316 (.ZN( u0_u3_n605 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U317 (.ZN( u0_u3_n530 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U318 (.ZN( u0_u3_n584 ) , .A1( u0_u3_n672 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U319 (.ZN( u0_u3_n444 ) , .A2( w3_28 ) , .A1( w3_29 ) );
  NOR4_X1 u0_u3_U32 (.A4( u0_u3_n529 ) , .A2( u0_u3_n530 ) , .A1( u0_u3_n531 ) , .ZN( u0_u3_n541 ) , .A3( u0_u3_n704 ) );
  NOR2_X1 u0_u3_U320 (.ZN( u0_u3_n468 ) , .A2( u0_u3_n849 ) , .A1( u0_u3_n850 ) );
  OAI222_X1 u0_u3_U321 (.B2( u0_u3_n750 ) , .B1( u0_u3_n751 ) , .A2( u0_u3_n752 ) , .ZN( u0_u3_n760 ) , .C2( u0_u3_n808 ) , .C1( u0_u3_n817 ) , .A1( u0_u3_n820 ) );
  INV_X1 u0_u3_U322 (.A( u0_u3_n789 ) , .ZN( u0_u3_n864 ) );
  NOR4_X1 u0_u3_U323 (.A4( u0_u3_n617 ) , .A3( u0_u3_n618 ) , .A1( u0_u3_n619 ) , .A2( u0_u3_n620 ) , .ZN( u0_u3_n621 ) );
  INV_X1 u0_u3_U324 (.ZN( u0_u3_n830 ) , .A( w3_25 ) );
  OAI22_X1 u0_u3_U325 (.B2( u0_u3_n753 ) , .B1( u0_u3_n754 ) , .A1( u0_u3_n755 ) , .ZN( u0_u3_n759 ) , .A2( u0_u3_n809 ) );
  OAI22_X1 u0_u3_U326 (.B2( u0_u3_n806 ) , .B1( u0_u3_n807 ) , .A2( u0_u3_n808 ) , .A1( u0_u3_n809 ) , .ZN( u0_u3_n811 ) );
  AOI21_X1 u0_u3_U327 (.ZN( u0_u3_n692 ) , .B2( u0_u3_n752 ) , .B1( u0_u3_n766 ) , .A( u0_u3_n809 ) );
  NAND2_X1 u0_u3_U328 (.A2( u0_u3_n765 ) , .A1( u0_u3_n809 ) , .ZN( u0_u3_n813 ) );
  NOR2_X1 u0_u3_U329 (.ZN( u0_u3_n573 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n809 ) );
  NOR4_X1 u0_u3_U33 (.A4( u0_u3_n535 ) , .A3( u0_u3_n536 ) , .A2( u0_u3_n537 ) , .ZN( u0_u3_n538 ) , .A1( u0_u3_n823 ) );
  NOR2_X1 u0_u3_U330 (.ZN( u0_u3_n614 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n809 ) );
  OAI22_X1 u0_u3_U331 (.ZN( u0_u3_n486 ) , .A1( u0_u3_n711 ) , .B2( u0_u3_n788 ) , .A2( u0_u3_n809 ) , .B1( u0_u3_n815 ) );
  AOI21_X1 u0_u3_U332 (.ZN( u0_u3_n480 ) , .A( u0_u3_n672 ) , .B1( u0_u3_n753 ) , .B2( u0_u3_n809 ) );
  INV_X1 u0_u3_U333 (.A( u0_u3_n809 ) , .ZN( u0_u3_n843 ) );
  OAI221_X1 u0_u3_U334 (.A( u0_u3_n786 ) , .C2( u0_u3_n787 ) , .B2( u0_u3_n788 ) , .B1( u0_u3_n789 ) , .ZN( u0_u3_n799 ) , .C1( u0_u3_n816 ) );
  NAND2_X1 u0_u3_U335 (.A1( u0_u3_n732 ) , .A2( u0_u3_n787 ) , .ZN( u0_u3_n814 ) );
  OAI22_X1 u0_u3_U336 (.ZN( u0_u3_n591 ) , .A2( u0_u3_n750 ) , .B2( u0_u3_n765 ) , .A1( u0_u3_n766 ) , .B1( u0_u3_n787 ) );
  AOI21_X1 u0_u3_U337 (.ZN( u0_u3_n595 ) , .B1( u0_u3_n731 ) , .B2( u0_u3_n787 ) , .A( u0_u3_n793 ) );
  NOR2_X1 u0_u3_U338 (.ZN( u0_u3_n807 ) , .A1( u0_u3_n856 ) , .A2( u0_u3_n863 ) );
  AOI21_X1 u0_u3_U339 (.ZN( u0_u3_n626 ) , .B1( u0_u3_n702 ) , .A( u0_u3_n782 ) , .B2( u0_u3_n787 ) );
  NOR4_X1 u0_u3_U34 (.A4( u0_u3_n532 ) , .A3( u0_u3_n533 ) , .ZN( u0_u3_n540 ) , .A2( u0_u3_n687 ) , .A1( u0_u3_n797 ) );
  NAND2_X2 u0_u3_U340 (.A1( u0_u3_n458 ) , .A2( u0_u3_n465 ) , .ZN( u0_u3_n753 ) );
  AOI222_X1 u0_u3_U341 (.ZN( u0_u3_n778 ) , .A1( u0_u3_n833 ) , .C1( u0_u3_n837 ) , .B2( u0_u3_n843 ) , .A2( u0_u3_n852 ) , .B1( u0_u3_n863 ) , .C2( u0_u3_n875 ) );
  AOI222_X1 u0_u3_U342 (.ZN( u0_u3_n609 ) , .A1( u0_u3_n833 ) , .C2( u0_u3_n839 ) , .B1( u0_u3_n844 ) , .A2( u0_u3_n858 ) , .B2( u0_u3_n863 ) , .C1( u0_u3_n870 ) );
  AOI21_X1 u0_u3_U343 (.ZN( u0_u3_n651 ) , .A( u0_u3_n765 ) , .B2( u0_u3_n787 ) , .B1( u0_u3_n795 ) );
  OAI22_X1 u0_u3_U344 (.ZN( u0_u3_n684 ) , .A1( u0_u3_n702 ) , .A2( u0_u3_n733 ) , .B2( u0_u3_n787 ) , .B1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U345 (.ZN( u0_u3_n654 ) , .A1( u0_u3_n787 ) , .A2( u0_u3_n791 ) );
  NOR2_X1 u0_u3_U346 (.ZN( u0_u3_n751 ) , .A1( u0_u3_n863 ) , .A2( u0_u3_n864 ) );
  NOR2_X1 u0_u3_U347 (.ZN( u0_u3_n455 ) , .A1( u0_u3_n860 ) , .A2( w3_30 ) );
  NOR2_X1 u0_u3_U348 (.ZN( u0_u3_n467 ) , .A2( w3_30 ) , .A1( w3_31 ) );
  AND2_X1 u0_u3_U349 (.ZN( u0_u3_n441 ) , .A2( u0_u3_n834 ) , .A1( u0_u3_n856 ) );
  NOR3_X1 u0_u3_U35 (.A3( u0_u3_n803 ) , .A2( u0_u3_n804 ) , .A1( u0_u3_n805 ) , .ZN( u0_u3_n828 ) );
  AND2_X1 u0_u3_U350 (.ZN( u0_u3_n442 ) , .A2( u0_u3_n845 ) , .A1( u0_u3_n863 ) );
  NOR3_X1 u0_u3_U351 (.A3( u0_u3_n441 ) , .A2( u0_u3_n442 ) , .A1( u0_u3_n579 ) , .ZN( u0_u3_n590 ) );
  INV_X1 u0_u3_U352 (.A( u0_u3_n815 ) , .ZN( u0_u3_n856 ) );
  INV_X1 u0_u3_U353 (.A( u0_u3_n787 ) , .ZN( u0_u3_n863 ) );
  INV_X1 u0_u3_U354 (.A( u0_u3_n806 ) , .ZN( u0_u3_n845 ) );
  INV_X1 u0_u3_U355 (.A( u0_u3_n41 ) , .ZN( u0_u3_n840 ) );
  NOR2_X1 u0_u3_U356 (.A1( u0_u3_n41 ) , .ZN( u0_u3_n773 ) , .A2( u0_u3_n818 ) );
  AOI21_X1 u0_u3_U357 (.B2( u0_u3_n41 ) , .ZN( u0_u3_n574 ) , .B1( u0_u3_n809 ) , .A( u0_u3_n815 ) );
  NOR2_X1 u0_u3_U358 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n665 ) , .A1( u0_u3_n732 ) );
  NOR2_X1 u0_u3_U359 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n635 ) , .A1( u0_u3_n727 ) );
  NAND4_X1 u0_u3_U36 (.A4( u0_u3_n660 ) , .A3( u0_u3_n661 ) , .A2( u0_u3_n662 ) , .A1( u0_u3_n663 ) , .ZN( u0_u3_n803 ) );
  NOR2_X1 u0_u3_U360 (.A2( u0_u3_n41 ) , .A1( u0_u3_n783 ) , .ZN( u0_u3_n823 ) );
  AOI21_X1 u0_u3_U361 (.B2( u0_u3_n41 ) , .ZN( u0_u3_n481 ) , .A( u0_u3_n752 ) , .B1( u0_u3_n782 ) );
  NOR2_X1 u0_u3_U362 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n569 ) , .A1( u0_u3_n766 ) );
  NOR2_X1 u0_u3_U363 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n719 ) , .A1( u0_u3_n795 ) );
  NOR2_X1 u0_u3_U364 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n597 ) , .A1( u0_u3_n731 ) );
  AOI21_X1 u0_u3_U365 (.A( u0_u3_n41 ) , .ZN( u0_u3_n555 ) , .B1( u0_u3_n672 ) , .B2( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U366 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n544 ) , .A1( u0_u3_n702 ) );
  NOR2_X1 u0_u3_U367 (.ZN( u0_u3_n583 ) , .A2( u0_u3_n700 ) , .A1( u0_u3_n794 ) );
  NOR4_X1 u0_u3_U368 (.A4( u0_u3_n779 ) , .A3( u0_u3_n780 ) , .A1( u0_u3_n781 ) , .ZN( u0_u3_n802 ) , .A2( u0_u3_n804 ) );
  NAND4_X1 u0_u3_U369 (.A4( u0_u3_n694 ) , .A3( u0_u3_n695 ) , .A1( u0_u3_n696 ) , .ZN( u0_u3_n779 ) , .A2( u0_u3_n874 ) );
  NOR3_X1 u0_u3_U37 (.A3( u0_u3_n654 ) , .A2( u0_u3_n655 ) , .A1( u0_u3_n656 ) , .ZN( u0_u3_n661 ) );
  AOI21_X1 u0_u3_U370 (.ZN( u0_u3_n596 ) , .B1( u0_u3_n753 ) , .A( u0_u3_n795 ) , .B2( u0_u3_n816 ) );
  AOI21_X1 u0_u3_U371 (.A( u0_u3_n815 ) , .B2( u0_u3_n816 ) , .B1( u0_u3_n817 ) , .ZN( u0_u3_n822 ) );
  OAI222_X1 u0_u3_U372 (.ZN( u0_u3_n508 ) , .C2( u0_u3_n628 ) , .B2( u0_u3_n650 ) , .B1( u0_u3_n750 ) , .A2( u0_u3_n751 ) , .C1( u0_u3_n808 ) , .A1( u0_u3_n809 ) );
  AOI21_X1 u0_u3_U373 (.B1( u0_u3_n628 ) , .ZN( u0_u3_n630 ) , .A( u0_u3_n766 ) , .B2( u0_u3_n817 ) );
  AOI21_X1 u0_u3_U374 (.ZN( u0_u3_n652 ) , .B1( u0_u3_n732 ) , .B2( u0_u3_n766 ) , .A( u0_u3_n816 ) );
  OAI21_X1 u0_u3_U375 (.A( u0_u3_n616 ) , .ZN( u0_u3_n619 ) , .B1( u0_u3_n628 ) , .B2( u0_u3_n787 ) );
  NOR2_X1 u0_u3_U376 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n769 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U377 (.A2( u0_u3_n816 ) , .A1( u0_u3_n818 ) , .ZN( u0_u3_n824 ) );
  NOR2_X1 u0_u3_U378 (.ZN( u0_u3_n581 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U379 (.A1( u0_u3_n439 ) , .ZN( u0_u3_n687 ) , .A2( u0_u3_n816 ) );
  NOR3_X1 u0_u3_U38 (.A3( u0_u3_n651 ) , .A2( u0_u3_n652 ) , .A1( u0_u3_n653 ) , .ZN( u0_u3_n662 ) );
  NOR2_X1 u0_u3_U380 (.ZN( u0_u3_n657 ) , .A1( u0_u3_n731 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U381 (.A1( u0_u3_n702 ) , .ZN( u0_u3_n771 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U382 (.ZN( u0_u3_n668 ) , .A1( u0_u3_n783 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U383 (.ZN( u0_u3_n634 ) , .A1( u0_u3_n727 ) , .A2( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U384 (.ZN( u0_u3_n475 ) , .A2( w3_26 ) , .A1( w3_27 ) );
  NOR2_X1 u0_u3_U385 (.ZN( u0_u3_n458 ) , .A1( u0_u3_n831 ) , .A2( w3_27 ) );
  INV_X1 u0_u3_U386 (.ZN( u0_u3_n832 ) , .A( w3_27 ) );
  NOR3_X1 u0_u3_U387 (.A3( u0_u3_n624 ) , .A2( u0_u3_n625 ) , .ZN( u0_u3_n639 ) , .A1( u0_u3_n728 ) );
  NOR4_X1 u0_u3_U388 (.A1( u0_u3_n587 ) , .ZN( u0_u3_n588 ) , .A3( u0_u3_n655 ) , .A2( u0_u3_n665 ) , .A4( u0_u3_n770 ) );
  OAI22_X1 u0_u3_U389 (.ZN( u0_u3_n640 ) , .A1( u0_u3_n702 ) , .B2( u0_u3_n731 ) , .A2( u0_u3_n765 ) , .B1( u0_u3_n819 ) );
  NOR3_X1 u0_u3_U39 (.A3( u0_u3_n657 ) , .A2( u0_u3_n658 ) , .A1( u0_u3_n659 ) , .ZN( u0_u3_n660 ) );
  AOI21_X1 u0_u3_U390 (.ZN( u0_u3_n502 ) , .B1( u0_u3_n683 ) , .A( u0_u3_n815 ) , .B2( u0_u3_n819 ) );
  OAI22_X1 u0_u3_U391 (.A1( u0_u3_n727 ) , .ZN( u0_u3_n729 ) , .B2( u0_u3_n753 ) , .B1( u0_u3_n815 ) , .A2( u0_u3_n819 ) );
  AOI21_X1 u0_u3_U392 (.A( u0_u3_n438 ) , .B2( u0_u3_n819 ) , .B1( u0_u3_n820 ) , .ZN( u0_u3_n821 ) );
  OAI22_X1 u0_u3_U393 (.A1( u0_u3_n438 ) , .ZN( u0_u3_n627 ) , .B1( u0_u3_n672 ) , .B2( u0_u3_n750 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U394 (.ZN( u0_u3_n522 ) , .A2( u0_u3_n702 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U395 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n691 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U396 (.A2( u0_u3_n439 ) , .ZN( u0_u3_n602 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U397 (.ZN( u0_u3_n534 ) , .A2( u0_u3_n783 ) , .A1( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U398 (.ZN( u0_u3_n561 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U399 (.ZN( u0_u3_n688 ) , .A1( u0_u3_n732 ) , .A2( u0_u3_n819 ) );
  NAND2_X1 u0_u3_U4 (.A1( u0_u3_n452 ) , .A2( u0_u3_n463 ) , .ZN( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U40 (.A4( u0_u3_n664 ) , .A3( u0_u3_n665 ) , .A2( u0_u3_n666 ) , .A1( u0_u3_n667 ) , .ZN( u0_u3_n680 ) );
  INV_X1 u0_u3_U400 (.A( u0_u3_n819 ) , .ZN( u0_u3_n834 ) );
  NAND2_X1 u0_u3_U401 (.ZN( u0_u3_n674 ) , .A1( u0_u3_n809 ) , .A2( u0_u3_n819 ) );
  NOR2_X1 u0_u3_U402 (.ZN( u0_u3_n465 ) , .A2( w3_24 ) , .A1( w3_25 ) );
  NOR2_X1 u0_u3_U403 (.ZN( u0_u3_n457 ) , .A1( u0_u3_n830 ) , .A2( w3_24 ) );
  INV_X1 u0_u3_U404 (.ZN( u0_u3_n829 ) , .A( w3_24 ) );
  INV_X1 u0_u3_U405 (.ZN( u0_u3_n850 ) , .A( w3_29 ) );
  NOR2_X1 u0_u3_U406 (.ZN( u0_u3_n451 ) , .A1( u0_u3_n849 ) , .A2( w3_29 ) );
  NAND4_X1 u0_u3_U407 (.ZN( u0_subword_3 ) , .A4( u0_u3_n707 ) , .A3( u0_u3_n708 ) , .A2( u0_u3_n709 ) , .A1( u0_u3_n710 ) );
  INV_X1 u0_u3_U408 (.A( u0_u3_n709 ) , .ZN( u0_u3_n878 ) );
  OAI22_X1 u0_u3_U409 (.B2( u0_u3_n747 ) , .ZN( u0_u3_n749 ) , .A2( u0_u3_n765 ) , .B1( u0_u3_n783 ) , .A1( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U41 (.A4( u0_u3_n668 ) , .A3( u0_u3_n669 ) , .A2( u0_u3_n670 ) , .A1( u0_u3_n671 ) , .ZN( u0_u3_n679 ) );
  OAI22_X1 u0_u3_U410 (.B1( u0_u3_n439 ) , .ZN( u0_u3_n499 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n783 ) , .B2( u0_u3_n809 ) );
  NOR2_X1 u0_u3_U411 (.ZN( u0_u3_n519 ) , .A1( u0_u3_n711 ) , .A2( u0_u3_n747 ) );
  OAI22_X1 u0_u3_U412 (.ZN( u0_u3_n713 ) , .A2( u0_u3_n731 ) , .B2( u0_u3_n732 ) , .A1( u0_u3_n747 ) , .B1( u0_u3_n816 ) );
  NOR2_X1 u0_u3_U413 (.A2( u0_u3_n747 ) , .ZN( u0_u3_n772 ) , .A1( u0_u3_n815 ) );
  OAI22_X1 u0_u3_U414 (.B1( u0_u3_n443 ) , .ZN( u0_u3_n447 ) , .A2( u0_u3_n731 ) , .A1( u0_u3_n747 ) , .B2( u0_u3_n752 ) );
  NOR2_X1 u0_u3_U415 (.ZN( u0_u3_n550 ) , .A1( u0_u3_n702 ) , .A2( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U416 (.ZN( u0_u3_n556 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n787 ) );
  NOR2_X1 u0_u3_U417 (.A2( u0_u3_n747 ) , .ZN( u0_u3_n758 ) , .A1( u0_u3_n808 ) );
  NOR2_X1 u0_u3_U418 (.A1( u0_u3_n672 ) , .ZN( u0_u3_n676 ) , .A2( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U419 (.ZN( u0_u3_n533 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n795 ) );
  NOR4_X1 u0_u3_U42 (.A3( u0_u3_n676 ) , .A1( u0_u3_n677 ) , .ZN( u0_u3_n678 ) , .A4( u0_u3_n718 ) , .A2( u0_u3_n861 ) );
  NOR2_X1 u0_u3_U420 (.ZN( u0_u3_n721 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n747 ) );
  NOR2_X1 u0_u3_U421 (.ZN( u0_u3_n585 ) , .A1( u0_u3_n747 ) , .A2( u0_u3_n818 ) );
  INV_X1 u0_u3_U422 (.A( u0_u3_n747 ) , .ZN( u0_u3_n839 ) );
  AOI21_X1 u0_u3_U423 (.ZN( u0_u3_n579 ) , .B2( u0_u3_n727 ) , .B1( u0_u3_n751 ) , .A( u0_u3_n788 ) );
  NAND4_X1 u0_u3_U424 (.A4( u0_u3_n636 ) , .A3( u0_u3_n637 ) , .A2( u0_u3_n638 ) , .A1( u0_u3_n639 ) , .ZN( u0_u3_n746 ) );
  INV_X1 u0_u3_U425 (.ZN( u0_u3_n851 ) , .A( w3_30 ) );
  INV_X1 u0_u3_U426 (.ZN( u0_u3_n860 ) , .A( w3_31 ) );
  NAND4_X1 u0_u3_U427 (.ZN( u0_subword_2 ) , .A4( u0_u3_n646 ) , .A3( u0_u3_n647 ) , .A2( u0_u3_n648 ) , .A1( u0_u3_n649 ) );
  AOI211_X1 u0_u3_U428 (.A( u0_u3_n640 ) , .ZN( u0_u3_n648 ) , .B( u0_u3_n746 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n856 ) );
  NOR2_X1 u0_u3_U429 (.A2( u0_u3_n41 ) , .ZN( u0_u3_n603 ) , .A1( u0_u3_n787 ) );
  NOR4_X1 u0_u3_U43 (.A1( u0_u3_n469 ) , .ZN( u0_u3_n470 ) , .A4( u0_u3_n545 ) , .A2( u0_u3_n557 ) , .A3( u0_u3_n617 ) );
  OAI222_X1 u0_u3_U430 (.A2( u0_u3_n672 ) , .ZN( u0_u3_n677 ) , .B1( u0_u3_n750 ) , .B2( u0_u3_n787 ) , .C2( u0_u3_n791 ) , .C1( u0_u3_n818 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U431 (.ZN( u0_u3_n613 ) , .A1( u0_u3_n787 ) , .A2( u0_u3_n819 ) );
  AOI21_X1 u0_u3_U432 (.A( u0_u3_n41 ) , .ZN( u0_u3_n503 ) , .B1( u0_u3_n711 ) , .B2( u0_u3_n789 ) );
  OAI22_X1 u0_u3_U433 (.ZN( u0_u3_n593 ) , .B1( u0_u3_n733 ) , .B2( u0_u3_n752 ) , .A2( u0_u3_n789 ) , .A1( u0_u3_n806 ) );
  NOR2_X1 u0_u3_U434 (.ZN( u0_u3_n656 ) , .A1( u0_u3_n765 ) , .A2( u0_u3_n789 ) );
  NAND2_X1 u0_u3_U435 (.A2( u0_u3_n752 ) , .A1( u0_u3_n789 ) , .ZN( u0_u3_n812 ) );
  NOR2_X1 u0_u3_U436 (.ZN( u0_u3_n557 ) , .A1( u0_u3_n789 ) , .A2( u0_u3_n816 ) );
  NAND3_X1 u0_u3_U437 (.ZN( u0_subword_6 ) , .A3( u0_u3_n800 ) , .A2( u0_u3_n801 ) , .A1( u0_u3_n802 ) );
  NAND3_X1 u0_u3_U438 (.ZN( u0_subword_5 ) , .A3( u0_u3_n761 ) , .A2( u0_u3_n762 ) , .A1( u0_u3_n763 ) );
  NAND3_X1 u0_u3_U439 (.ZN( u0_subword_4 ) , .A3( u0_u3_n741 ) , .A2( u0_u3_n742 ) , .A1( u0_u3_n743 ) );
  AOI221_X1 u0_u3_U44 (.ZN( u0_u3_n471 ) , .C2( u0_u3_n717 ) , .B2( u0_u3_n834 ) , .C1( u0_u3_n847 ) , .B1( u0_u3_n862 ) , .A( u0_u3_n866 ) );
  NAND3_X1 u0_u3_U440 (.A3( u0_u3_n678 ) , .A2( u0_u3_n679 ) , .A1( u0_u3_n680 ) , .ZN( u0_u3_n810 ) );
  NAND3_X1 u0_u3_U441 (.ZN( u0_u3_n641 ) , .A3( u0_u3_n711 ) , .A2( u0_u3_n727 ) , .A1( u0_u3_n795 ) );
  NAND3_X1 u0_u3_U442 (.A3( u0_u3_n621 ) , .A2( u0_u3_n622 ) , .A1( u0_u3_n623 ) , .ZN( u0_u3_n728 ) );
  NAND3_X1 u0_u3_U443 (.A3( u0_u3_n588 ) , .A2( u0_u3_n589 ) , .A1( u0_u3_n590 ) , .ZN( u0_u3_n624 ) );
  NAND3_X1 u0_u3_U444 (.ZN( u0_u3_n568 ) , .A3( u0_u3_n683 ) , .A2( u0_u3_n753 ) , .A1( u0_u3_n788 ) );
  NAND3_X1 u0_u3_U445 (.A3( u0_u3_n526 ) , .A2( u0_u3_n527 ) , .A1( u0_u3_n528 ) , .ZN( u0_u3_n745 ) );
  NAND3_X1 u0_u3_U446 (.A3( u0_u3_n515 ) , .A1( u0_u3_n516 ) , .ZN( u0_u3_n611 ) , .A2( u0_u3_n873 ) );
  NAND3_X1 u0_u3_U447 (.A3( u0_u3_n470 ) , .A2( u0_u3_n471 ) , .A1( u0_u3_n472 ) , .ZN( u0_u3_n780 ) );
  NOR2_X1 u0_u3_U448 (.ZN( u0_u3_n615 ) , .A1( u0_u3_n782 ) , .A2( u0_u3_n789 ) );
  NOR2_X1 u0_u3_U449 (.ZN( u0_u3_n720 ) , .A2( u0_u3_n747 ) , .A1( u0_u3_n789 ) );
  NOR4_X1 u0_u3_U45 (.A4( u0_u3_n517 ) , .A3( u0_u3_n518 ) , .A2( u0_u3_n519 ) , .A1( u0_u3_n520 ) , .ZN( u0_u3_n527 ) );
  NOR2_X1 u0_u3_U450 (.ZN( u0_u3_n704 ) , .A2( u0_u3_n789 ) , .A1( u0_u3_n820 ) );
  NOR2_X1 u0_u3_U451 (.A1( u0_u3_n733 ) , .ZN( u0_u3_n768 ) , .A2( u0_u3_n789 ) );
  INV_X1 u0_u3_U452 (.ZN( u0_u3_n849 ) , .A( w3_28 ) );
  NOR4_X1 u0_u3_U46 (.A3( u0_u3_n524 ) , .A1( u0_u3_n525 ) , .ZN( u0_u3_n526 ) , .A2( u0_u3_n676 ) , .A4( u0_u3_n772 ) );
  NAND4_X1 u0_u3_U47 (.A4( u0_u3_n576 ) , .A3( u0_u3_n577 ) , .A1( u0_u3_n578 ) , .ZN( u0_u3_n726 ) , .A2( u0_u3_n876 ) );
  NOR4_X1 u0_u3_U48 (.A4( u0_u3_n572 ) , .A3( u0_u3_n573 ) , .A2( u0_u3_n574 ) , .A1( u0_u3_n575 ) , .ZN( u0_u3_n576 ) );
  INV_X1 u0_u3_U49 (.A( u0_u3_n610 ) , .ZN( u0_u3_n876 ) );
  NAND2_X1 u0_u3_U5 (.A1( u0_u3_n456 ) , .A2( u0_u3_n475 ) , .ZN( u0_u3_n788 ) );
  NAND4_X1 u0_u3_U50 (.A4( u0_u3_n459 ) , .A3( u0_u3_n460 ) , .A2( u0_u3_n461 ) , .A1( u0_u3_n462 ) , .ZN( u0_u3_n682 ) );
  NOR3_X1 u0_u3_U51 (.ZN( u0_u3_n460 ) , .A3( u0_u3_n533 ) , .A1( u0_u3_n558 ) , .A2( u0_u3_n573 ) );
  NOR4_X1 u0_u3_U52 (.ZN( u0_u3_n459 ) , .A2( u0_u3_n520 ) , .A1( u0_u3_n546 ) , .A3( u0_u3_n582 ) , .A4( u0_u3_n618 ) );
  NOR4_X1 u0_u3_U53 (.ZN( u0_u3_n461 ) , .A2( u0_u3_n512 ) , .A1( u0_u3_n602 ) , .A4( u0_u3_n631 ) , .A3( u0_u3_n714 ) );
  NAND4_X1 u0_u3_U54 (.A4( u0_u3_n722 ) , .A3( u0_u3_n723 ) , .A2( u0_u3_n724 ) , .ZN( u0_u3_n744 ) , .A1( u0_u3_n859 ) );
  INV_X1 u0_u3_U55 (.A( u0_u3_n712 ) , .ZN( u0_u3_n859 ) );
  NOR4_X1 u0_u3_U56 (.A4( u0_u3_n718 ) , .A3( u0_u3_n719 ) , .A2( u0_u3_n720 ) , .A1( u0_u3_n721 ) , .ZN( u0_u3_n722 ) );
  NOR3_X1 u0_u3_U57 (.ZN( u0_u3_n483 ) , .A2( u0_u3_n511 ) , .A3( u0_u3_n604 ) , .A1( u0_u3_n613 ) );
  NOR4_X1 u0_u3_U58 (.ZN( u0_u3_n484 ) , .A3( u0_u3_n535 ) , .A4( u0_u3_n548 ) , .A2( u0_u3_n570 ) , .A1( u0_u3_n720 ) );
  AOI211_X1 u0_u3_U59 (.B( u0_u3_n480 ) , .A( u0_u3_n481 ) , .ZN( u0_u3_n485 ) , .C2( u0_u3_n836 ) , .C1( u0_u3_n863 ) );
  NOR3_X1 u0_u3_U6 (.ZN( u0_u3_n601 ) , .A1( u0_u3_n611 ) , .A3( u0_u3_n726 ) , .A2( u0_u3_n745 ) );
  INV_X1 u0_u3_U60 (.A( u0_u3_n682 ) , .ZN( u0_u3_n874 ) );
  NOR4_X1 u0_u3_U61 (.A4( u0_u3_n690 ) , .A3( u0_u3_n691 ) , .A2( u0_u3_n692 ) , .A1( u0_u3_n693 ) , .ZN( u0_u3_n694 ) );
  AOI221_X1 u0_u3_U62 (.A( u0_u3_n684 ) , .ZN( u0_u3_n695 ) , .B2( u0_u3_n842 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n864 ) , .B1( u0_u3_n867 ) );
  NAND4_X1 u0_u3_U63 (.A4( u0_u3_n476 ) , .A3( u0_u3_n477 ) , .A2( u0_u3_n478 ) , .A1( u0_u3_n479 ) , .ZN( u0_u3_n681 ) );
  NOR4_X1 u0_u3_U64 (.A4( u0_u3_n473 ) , .ZN( u0_u3_n479 ) , .A3( u0_u3_n559 ) , .A1( u0_u3_n738 ) , .A2( u0_u3_n758 ) );
  NOR4_X1 u0_u3_U65 (.ZN( u0_u3_n477 ) , .A1( u0_u3_n509 ) , .A3( u0_u3_n547 ) , .A2( u0_u3_n586 ) , .A4( u0_u3_n719 ) );
  NOR4_X1 u0_u3_U66 (.ZN( u0_u3_n476 ) , .A2( u0_u3_n524 ) , .A4( u0_u3_n597 ) , .A1( u0_u3_n612 ) , .A3( u0_u3_n632 ) );
  NAND4_X1 u0_u3_U67 (.A4( u0_u3_n551 ) , .A3( u0_u3_n552 ) , .A2( u0_u3_n553 ) , .A1( u0_u3_n554 ) , .ZN( u0_u3_n748 ) );
  AOI211_X1 u0_u3_U68 (.B( u0_u3_n542 ) , .A( u0_u3_n543 ) , .ZN( u0_u3_n554 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n853 ) );
  NOR3_X1 u0_u3_U69 (.ZN( u0_u3_n552 ) , .A2( u0_u3_n654 ) , .A1( u0_u3_n670 ) , .A3( u0_u3_n774 ) );
  NOR3_X1 u0_u3_U7 (.ZN( u0_u3_n507 ) , .A2( u0_u3_n682 ) , .A3( u0_u3_n780 ) , .A1( u0_u3_n878 ) );
  NOR4_X1 u0_u3_U70 (.A4( u0_u3_n544 ) , .A3( u0_u3_n545 ) , .A2( u0_u3_n546 ) , .ZN( u0_u3_n553 ) , .A1( u0_u3_n691 ) );
  NOR4_X1 u0_u3_U71 (.A4( u0_u3_n612 ) , .A3( u0_u3_n613 ) , .A2( u0_u3_n614 ) , .A1( u0_u3_n615 ) , .ZN( u0_u3_n622 ) );
  NOR4_X1 u0_u3_U72 (.ZN( u0_u3_n623 ) , .A1( u0_u3_n659 ) , .A3( u0_u3_n669 ) , .A4( u0_u3_n685 ) , .A2( u0_u3_n769 ) );
  INV_X1 u0_u3_U73 (.A( u0_u3_n765 ) , .ZN( u0_u3_n833 ) );
  NOR2_X1 u0_u3_U74 (.ZN( u0_u3_n650 ) , .A1( u0_u3_n856 ) , .A2( u0_u3_n870 ) );
  NOR4_X1 u0_u3_U75 (.A4( u0_u3_n580 ) , .A3( u0_u3_n581 ) , .A2( u0_u3_n582 ) , .ZN( u0_u3_n589 ) , .A1( u0_u3_n686 ) );
  INV_X1 u0_u3_U76 (.A( u0_u3_n818 ) , .ZN( u0_u3_n857 ) );
  OR4_X1 u0_u3_U77 (.A4( u0_u3_n685 ) , .A3( u0_u3_n686 ) , .A2( u0_u3_n687 ) , .A1( u0_u3_n688 ) , .ZN( u0_u3_n693 ) );
  OR4_X1 u0_u3_U78 (.ZN( u0_u3_n469 ) , .A4( u0_u3_n521 ) , .A3( u0_u3_n532 ) , .A2( u0_u3_n581 ) , .A1( u0_u3_n715 ) );
  OR4_X1 u0_u3_U79 (.A4( u0_u3_n569 ) , .A3( u0_u3_n570 ) , .A2( u0_u3_n571 ) , .ZN( u0_u3_n575 ) , .A1( u0_u3_n668 ) );
  NOR3_X1 u0_u3_U8 (.A2( u0_u3_n610 ) , .A1( u0_u3_n611 ) , .ZN( u0_u3_n649 ) , .A3( u0_u3_n725 ) );
  OR4_X1 u0_u3_U80 (.A4( u0_u3_n521 ) , .A2( u0_u3_n522 ) , .A1( u0_u3_n523 ) , .ZN( u0_u3_n525 ) , .A3( u0_u3_n824 ) );
  OR4_X1 u0_u3_U81 (.A4( u0_u3_n583 ) , .A3( u0_u3_n584 ) , .A2( u0_u3_n585 ) , .A1( u0_u3_n586 ) , .ZN( u0_u3_n587 ) );
  OR4_X1 u0_u3_U82 (.ZN( u0_u3_n495 ) , .A4( u0_u3_n537 ) , .A2( u0_u3_n550 ) , .A1( u0_u3_n562 ) , .A3( u0_u3_n635 ) );
  NOR4_X1 u0_u3_U83 (.A4( u0_u3_n512 ) , .A2( u0_u3_n513 ) , .A1( u0_u3_n514 ) , .ZN( u0_u3_n515 ) , .A3( u0_u3_n673 ) );
  INV_X1 u0_u3_U84 (.A( u0_u3_n508 ) , .ZN( u0_u3_n873 ) );
  OR3_X1 u0_u3_U85 (.A3( u0_u3_n509 ) , .A2( u0_u3_n510 ) , .A1( u0_u3_n511 ) , .ZN( u0_u3_n514 ) );
  INV_X1 u0_u3_U86 (.A( u0_u3_n757 ) , .ZN( u0_u3_n871 ) );
  AOI221_X1 u0_u3_U87 (.A( u0_u3_n716 ) , .B2( u0_u3_n717 ) , .ZN( u0_u3_n723 ) , .C1( u0_u3_n835 ) , .B1( u0_u3_n841 ) , .C2( u0_u3_n865 ) );
  OR2_X1 u0_u3_U88 (.A2( u0_u3_n714 ) , .A1( u0_u3_n715 ) , .ZN( u0_u3_n716 ) );
  INV_X1 u0_u3_U89 (.A( u0_u3_n466 ) , .ZN( u0_u3_n866 ) );
  NOR3_X1 u0_u3_U9 (.A3( u0_u3_n725 ) , .A1( u0_u3_n726 ) , .ZN( u0_u3_n743 ) , .A2( u0_u3_n744 ) );
  NAND2_X1 u0_u3_U90 (.A1( u0_u3_n454 ) , .A2( u0_u3_n456 ) , .ZN( u0_u3_n765 ) );
  AOI22_X1 u0_u3_U91 (.ZN( u0_u3_n699 ) , .A1( u0_u3_n833 ) , .B2( u0_u3_n845 ) , .A2( u0_u3_n867 ) , .B1( u0_u3_n870 ) );
  NOR3_X1 u0_u3_U92 (.ZN( u0_u3_n755 ) , .A2( u0_u3_n855 ) , .A1( u0_u3_n865 ) , .A3( u0_u3_n867 ) );
  NOR2_X1 u0_u3_U93 (.ZN( u0_u3_n754 ) , .A2( u0_u3_n854 ) , .A1( u0_u3_n862 ) );
  AOI211_X1 u0_u3_U94 (.A( u0_u3_n499 ) , .ZN( u0_u3_n506 ) , .B( u0_u3_n805 ) , .C2( u0_u3_n841 ) , .C1( u0_u3_n853 ) );
  AOI211_X1 u0_u3_U95 (.B( u0_u3_n810 ) , .A( u0_u3_n811 ) , .ZN( u0_u3_n827 ) , .C1( u0_u3_n844 ) , .C2( u0_u3_n852 ) );
  NAND2_X1 u0_u3_U96 (.A1( u0_u3_n450 ) , .A2( u0_u3_n468 ) , .ZN( u0_u3_n752 ) );
  INV_X1 u0_u3_U97 (.A( u0_u3_n733 ) , .ZN( u0_u3_n841 ) );
  AOI221_X1 u0_u3_U98 (.B2( u0_u3_n440 ) , .A( u0_u3_n492 ) , .ZN( u0_u3_n497 ) , .C2( u0_u3_n843 ) , .C1( u0_u3_n853 ) , .B1( u0_u3_n862 ) );
  INV_X1 u0_u3_U99 (.A( u0_u3_n781 ) , .ZN( u0_u3_n869 ) );
  NOR2_X1 us01_U10 (.ZN( us01_n573 ) , .A1( us01_n620 ) , .A2( us01_n743 ) );
  AOI211_X1 us01_U100 (.B( us01_n537 ) , .A( us01_n538 ) , .ZN( us01_n549 ) , .C2( us01_n837 ) , .C1( us01_n849 ) );
  NOR4_X1 us01_U101 (.A4( us01_n542 ) , .A3( us01_n543 ) , .A2( us01_n544 ) , .A1( us01_n545 ) , .ZN( us01_n546 ) );
  NOR4_X1 us01_U102 (.A4( us01_n607 ) , .A3( us01_n608 ) , .A2( us01_n609 ) , .A1( us01_n610 ) , .ZN( us01_n617 ) );
  NOR4_X1 us01_U103 (.ZN( us01_n618 ) , .A1( us01_n654 ) , .A3( us01_n664 ) , .A4( us01_n680 ) , .A2( us01_n764 ) );
  NOR4_X1 us01_U104 (.A4( us01_n612 ) , .A3( us01_n613 ) , .A2( us01_n614 ) , .A1( us01_n615 ) , .ZN( us01_n616 ) );
  NOR2_X1 us01_U105 (.ZN( us01_n684 ) , .A1( us01_n829 ) , .A2( us01_n830 ) );
  NAND4_X1 us01_U106 (.A4( us01_n471 ) , .A3( us01_n472 ) , .A2( us01_n473 ) , .A1( us01_n474 ) , .ZN( us01_n676 ) );
  NOR4_X1 us01_U107 (.A4( us01_n468 ) , .ZN( us01_n474 ) , .A3( us01_n554 ) , .A1( us01_n733 ) , .A2( us01_n753 ) );
  NOR4_X1 us01_U108 (.ZN( us01_n473 ) , .A1( us01_n529 ) , .A3( us01_n566 ) , .A4( us01_n598 ) , .A2( us01_n640 ) );
  NOR4_X1 us01_U109 (.ZN( us01_n472 ) , .A1( us01_n504 ) , .A3( us01_n542 ) , .A2( us01_n581 ) , .A4( us01_n714 ) );
  NOR2_X1 us01_U11 (.ZN( us01_n493 ) , .A1( us01_n676 ) , .A2( us01_n692 ) );
  NAND4_X1 us01_U110 (.A4( us01_n689 ) , .A3( us01_n690 ) , .A1( us01_n691 ) , .ZN( us01_n774 ) , .A2( us01_n870 ) );
  INV_X1 us01_U111 (.A( us01_n677 ) , .ZN( us01_n870 ) );
  AOI221_X1 us01_U112 (.A( us01_n679 ) , .ZN( us01_n690 ) , .B2( us01_n838 ) , .C1( us01_n840 ) , .C2( us01_n860 ) , .B1( us01_n863 ) );
  NOR4_X1 us01_U113 (.A4( us01_n685 ) , .A3( us01_n686 ) , .A2( us01_n687 ) , .A1( us01_n688 ) , .ZN( us01_n689 ) );
  NOR2_X1 us01_U114 (.ZN( us01_n731 ) , .A2( us01_n830 ) , .A1( us01_n843 ) );
  NAND4_X1 us01_U115 (.A4( us01_n717 ) , .A3( us01_n718 ) , .A2( us01_n719 ) , .ZN( us01_n739 ) , .A1( us01_n855 ) );
  AOI221_X1 us01_U116 (.A( us01_n708 ) , .ZN( us01_n719 ) , .C2( us01_n842 ) , .B2( us01_n843 ) , .C1( us01_n859 ) , .B1( us01_n860 ) );
  INV_X1 us01_U117 (.A( us01_n707 ) , .ZN( us01_n855 ) );
  NOR4_X1 us01_U118 (.A4( us01_n713 ) , .A3( us01_n714 ) , .A2( us01_n715 ) , .A1( us01_n716 ) , .ZN( us01_n717 ) );
  NOR2_X1 us01_U119 (.ZN( us01_n645 ) , .A1( us01_n852 ) , .A2( us01_n866 ) );
  NOR2_X1 us01_U12 (.A1( us01_n676 ) , .ZN( us01_n691 ) , .A2( us01_n805 ) );
  NAND4_X1 us01_U120 (.A4( us01_n571 ) , .A3( us01_n572 ) , .A1( us01_n573 ) , .ZN( us01_n721 ) , .A2( us01_n872 ) );
  AOI221_X1 us01_U121 (.A( us01_n562 ) , .C2( us01_n563 ) , .ZN( us01_n572 ) , .B2( us01_n843 ) , .B1( us01_n850 ) , .C1( us01_n851 ) );
  NOR4_X1 us01_U122 (.A4( us01_n567 ) , .A3( us01_n568 ) , .A2( us01_n569 ) , .A1( us01_n570 ) , .ZN( us01_n571 ) );
  INV_X1 us01_U123 (.A( us01_n605 ) , .ZN( us01_n872 ) );
  NAND4_X1 us01_U124 (.A4( us01_n491 ) , .A3( us01_n492 ) , .A1( us01_n493 ) , .ZN( us01_n800 ) , .A2( us01_n865 ) );
  AOI221_X1 us01_U125 (.A( us01_n487 ) , .ZN( us01_n492 ) , .B2( us01_n834 ) , .C2( us01_n839 ) , .C1( us01_n849 ) , .B1( us01_n858 ) );
  INV_X1 us01_U126 (.A( us01_n776 ) , .ZN( us01_n865 ) );
  NOR4_X1 us01_U127 (.A2( us01_n489 ) , .A1( us01_n490 ) , .ZN( us01_n491 ) , .A3( us01_n578 ) , .A4( us01_n610 ) );
  NOR4_X1 us01_U128 (.A3( us01_n753 ) , .A2( us01_n754 ) , .A1( us01_n755 ) , .ZN( us01_n756 ) , .A4( us01_n867 ) );
  AOI211_X1 us01_U129 (.B( us01_n743 ) , .A( us01_n744 ) , .ZN( us01_n757 ) , .C1( us01_n830 ) , .C2( us01_n851 ) );
  NOR3_X1 us01_U13 (.ZN( us01_n502 ) , .A2( us01_n677 ) , .A3( us01_n775 ) , .A1( us01_n874 ) );
  NOR3_X1 us01_U130 (.A3( us01_n739 ) , .A2( us01_n740 ) , .A1( us01_n741 ) , .ZN( us01_n758 ) );
  NOR4_X1 us01_U131 (.A4( us01_n732 ) , .A3( us01_n733 ) , .A2( us01_n734 ) , .A1( us01_n735 ) , .ZN( us01_n736 ) );
  AOI211_X1 us01_U132 (.B( us01_n723 ) , .A( us01_n724 ) , .ZN( us01_n737 ) , .C1( us01_n841 ) , .C2( us01_n853 ) );
  NOR3_X1 us01_U133 (.A3( us01_n720 ) , .A1( us01_n721 ) , .ZN( us01_n738 ) , .A2( us01_n739 ) );
  INV_X1 us01_U134 (.A( us01_n760 ) , .ZN( us01_n828 ) );
  NAND4_X1 us01_U135 (.ZN( sa01_sr_3 ) , .A4( us01_n702 ) , .A3( us01_n703 ) , .A2( us01_n704 ) , .A1( us01_n705 ) );
  NOR4_X1 us01_U136 (.A4( us01_n698 ) , .A3( us01_n699 ) , .A2( us01_n700 ) , .A1( us01_n701 ) , .ZN( us01_n702 ) );
  AOI211_X1 us01_U137 (.B( us01_n692 ) , .A( us01_n693 ) , .ZN( us01_n703 ) , .C2( us01_n829 ) , .C1( us01_n849 ) );
  NOR2_X1 us01_U138 (.ZN( us01_n705 ) , .A2( us01_n774 ) , .A1( us01_n798 ) );
  OR4_X1 us01_U139 (.A4( us01_n680 ) , .A3( us01_n681 ) , .A2( us01_n682 ) , .A1( us01_n683 ) , .ZN( us01_n688 ) );
  INV_X1 us01_U14 (.A( us01_n704 ) , .ZN( us01_n874 ) );
  OR4_X1 us01_U140 (.ZN( us01_n464 ) , .A4( us01_n516 ) , .A3( us01_n527 ) , .A2( us01_n576 ) , .A1( us01_n710 ) );
  OR4_X1 us01_U141 (.A4( us01_n564 ) , .A3( us01_n565 ) , .A2( us01_n566 ) , .ZN( us01_n570 ) , .A1( us01_n663 ) );
  OR4_X1 us01_U142 (.A4( us01_n516 ) , .A2( us01_n517 ) , .A1( us01_n518 ) , .ZN( us01_n520 ) , .A3( us01_n819 ) );
  OR4_X1 us01_U143 (.ZN( us01_n490 ) , .A4( us01_n532 ) , .A2( us01_n545 ) , .A1( us01_n557 ) , .A3( us01_n630 ) );
  OR4_X1 us01_U144 (.A4( us01_n578 ) , .A3( us01_n579 ) , .A2( us01_n580 ) , .A1( us01_n581 ) , .ZN( us01_n582 ) );
  INV_X1 us01_U145 (.A( us01_n695 ) , .ZN( us01_n836 ) );
  NAND2_X1 us01_U146 (.ZN( us01_n611 ) , .A2( us01_n835 ) , .A1( us01_n871 ) );
  OR3_X1 us01_U147 (.A3( us01_n504 ) , .A2( us01_n505 ) , .A1( us01_n506 ) , .ZN( us01_n509 ) );
  AOI221_X1 us01_U148 (.A( us01_n711 ) , .B2( us01_n712 ) , .ZN( us01_n718 ) , .C1( us01_n830 ) , .B1( us01_n837 ) , .C2( us01_n861 ) );
  OR2_X1 us01_U149 (.A2( us01_n709 ) , .A1( us01_n710 ) , .ZN( us01_n711 ) );
  INV_X1 us01_U15 (.A( us01_n678 ) , .ZN( us01_n838 ) );
  INV_X1 us01_U150 (.A( us01_n461 ) , .ZN( us01_n862 ) );
  OAI21_X1 us01_U151 (.ZN( us01_n461 ) , .B1( us01_n807 ) , .A( us01_n832 ) , .B2( us01_n849 ) );
  INV_X1 us01_U152 (.A( us01_n752 ) , .ZN( us01_n867 ) );
  OAI21_X1 us01_U153 (.B1( us01_n751 ) , .ZN( us01_n752 ) , .A( us01_n843 ) , .B2( us01_n866 ) );
  INV_X1 us01_U154 (.A( us01_n670 ) , .ZN( us01_n857 ) );
  AOI21_X1 us01_U155 (.A( us01_n668 ) , .B1( us01_n669 ) , .ZN( us01_n670 ) , .B2( us01_n854 ) );
  AOI222_X1 us01_U156 (.ZN( us01_n658 ) , .A2( us01_n837 ) , .B1( us01_n839 ) , .C2( us01_n843 ) , .A1( us01_n858 ) , .C1( us01_n861 ) , .B2( us01_n868 ) );
  INV_X1 us01_U157 (.A( us01_n645 ) , .ZN( us01_n868 ) );
  OAI22_X1 us01_U158 (.ZN( us01_n481 ) , .A1( us01_n706 ) , .B2( us01_n783 ) , .A2( us01_n804 ) , .B1( us01_n810 ) );
  OAI22_X1 us01_U159 (.ZN( us01_n635 ) , .A1( us01_n697 ) , .B2( us01_n726 ) , .A2( us01_n760 ) , .B1( us01_n814 ) );
  NOR4_X1 us01_U16 (.A4( us01_n443 ) , .A3( us01_n444 ) , .A2( us01_n514 ) , .A1( us01_n539 ) , .ZN( us01_n704 ) );
  OAI222_X1 us01_U160 (.ZN( us01_n503 ) , .C2( us01_n623 ) , .B2( us01_n645 ) , .B1( us01_n745 ) , .A2( us01_n746 ) , .C1( us01_n803 ) , .A1( us01_n804 ) );
  OAI222_X1 us01_U161 (.B2( us01_n745 ) , .B1( us01_n746 ) , .A2( us01_n747 ) , .ZN( us01_n755 ) , .C2( us01_n803 ) , .C1( us01_n812 ) , .A1( us01_n815 ) );
  OAI222_X1 us01_U162 (.B2( us01_n706 ) , .ZN( us01_n707 ) , .C2( us01_n722 ) , .B1( us01_n745 ) , .A1( us01_n804 ) , .C1( us01_n812 ) , .A2( us01_n813 ) );
  AOI22_X1 us01_U163 (.ZN( us01_n694 ) , .A1( us01_n828 ) , .B2( us01_n841 ) , .A2( us01_n863 ) , .B1( us01_n866 ) );
  AOI22_X1 us01_U164 (.A2( us01_n780 ) , .ZN( us01_n781 ) , .B2( us01_n829 ) , .A1( us01_n832 ) , .B1( us01_n861 ) );
  INV_X1 us01_U165 (.A( us01_n728 ) , .ZN( us01_n837 ) );
  AOI221_X1 us01_U166 (.A( us01_n762 ) , .ZN( us01_n772 ) , .C2( us01_n808 ) , .B2( us01_n833 ) , .C1( us01_n853 ) , .B1( us01_n864 ) );
  AOI21_X1 us01_U167 (.B2( us01_n761 ) , .ZN( us01_n762 ) , .A( us01_n786 ) , .B1( us01_n790 ) );
  INV_X1 us01_U168 (.A( us01_n759 ) , .ZN( us01_n833 ) );
  INV_X1 us01_U169 (.A( us01_n788 ) , .ZN( us01_n830 ) );
  OR3_X1 us01_U17 (.ZN( us01_n444 ) , .A1( us01_n526 ) , .A3( us01_n575 ) , .A2( us01_n873 ) );
  OAI221_X1 us01_U170 (.A( us01_n725 ) , .C2( us01_n726 ) , .B2( us01_n727 ) , .B1( us01_n728 ) , .ZN( us01_n735 ) , .C1( us01_n815 ) );
  AOI22_X1 us01_U171 (.ZN( us01_n725 ) , .B1( us01_n830 ) , .A2( us01_n836 ) , .A1( us01_n861 ) , .B2( us01_n864 ) );
  NAND2_X1 us01_U172 (.A1( us01_n449 ) , .A2( us01_n451 ) , .ZN( us01_n760 ) );
  OAI22_X1 us01_U173 (.ZN( us01_n622 ) , .B1( us01_n667 ) , .B2( us01_n745 ) , .A1( us01_n813 ) , .A2( us01_n814 ) );
  OAI22_X1 us01_U174 (.A1( us01_n722 ) , .ZN( us01_n724 ) , .B2( us01_n748 ) , .B1( us01_n810 ) , .A2( us01_n814 ) );
  OAI22_X1 us01_U175 (.ZN( us01_n487 ) , .A1( us01_n722 ) , .B2( us01_n726 ) , .B1( us01_n728 ) , .A2( us01_n777 ) );
  OAI22_X1 us01_U176 (.B2( us01_n777 ) , .B1( us01_n778 ) , .ZN( us01_n779 ) , .A2( us01_n812 ) , .A1( us01_n813 ) );
  OAI22_X1 us01_U177 (.B2( us01_n748 ) , .B1( us01_n749 ) , .A1( us01_n750 ) , .ZN( us01_n754 ) , .A2( us01_n804 ) );
  NOR3_X1 us01_U178 (.ZN( us01_n750 ) , .A2( us01_n851 ) , .A1( us01_n861 ) , .A3( us01_n863 ) );
  NOR2_X1 us01_U179 (.ZN( us01_n749 ) , .A2( us01_n850 ) , .A1( us01_n858 ) );
  OR4_X1 us01_U18 (.A4( us01_n440 ) , .A2( us01_n441 ) , .A1( us01_n442 ) , .ZN( us01_n443 ) , .A3( us01_n551 ) );
  INV_X1 us01_U180 (.A( us01_n803 ) , .ZN( us01_n858 ) );
  OAI22_X1 us01_U181 (.B2( us01_n742 ) , .ZN( us01_n744 ) , .A2( us01_n760 ) , .B1( us01_n778 ) , .A1( us01_n790 ) );
  OAI22_X1 us01_U182 (.ZN( us01_n494 ) , .A2( us01_n742 ) , .A1( us01_n778 ) , .B1( us01_n789 ) , .B2( us01_n804 ) );
  OAI22_X1 us01_U183 (.B2( us01_n801 ) , .B1( us01_n802 ) , .A2( us01_n803 ) , .A1( us01_n804 ) , .ZN( us01_n806 ) );
  OAI22_X1 us01_U184 (.ZN( us01_n693 ) , .A2( us01_n728 ) , .A1( us01_n778 ) , .B1( us01_n789 ) , .B2( us01_n815 ) );
  NOR2_X1 us01_U185 (.ZN( us01_n713 ) , .A1( us01_n803 ) , .A2( us01_n815 ) );
  NOR2_X1 us01_U186 (.A1( us01_n697 ) , .ZN( us01_n766 ) , .A2( us01_n811 ) );
  INV_X1 us01_U187 (.A( us01_n786 ) , .ZN( us01_n843 ) );
  NOR2_X1 us01_U188 (.ZN( us01_n539 ) , .A2( us01_n695 ) , .A1( us01_n697 ) );
  INV_X1 us01_U189 (.A( us01_n742 ) , .ZN( us01_n835 ) );
  INV_X1 us01_U19 (.A( us01_n611 ) , .ZN( us01_n873 ) );
  INV_X1 us01_U190 (.A( us01_n814 ) , .ZN( us01_n829 ) );
  INV_X1 us01_U191 (.A( us01_n812 ) , .ZN( us01_n831 ) );
  OAI22_X1 us01_U192 (.B1( us01_n488 ) , .ZN( us01_n489 ) , .A1( us01_n684 ) , .A2( us01_n761 ) , .B2( us01_n815 ) );
  NOR3_X1 us01_U193 (.ZN( us01_n488 ) , .A1( us01_n780 ) , .A2( us01_n848 ) , .A3( us01_n861 ) );
  NOR2_X1 us01_U194 (.A2( us01_n742 ) , .ZN( us01_n753 ) , .A1( us01_n803 ) );
  NOR2_X1 us01_U195 (.ZN( us01_n733 ) , .A2( us01_n801 ) , .A1( us01_n803 ) );
  INV_X1 us01_U196 (.A( us01_n790 ) , .ZN( us01_n849 ) );
  NOR2_X1 us01_U197 (.A2( us01_n742 ) , .ZN( us01_n767 ) , .A1( us01_n810 ) );
  NOR2_X1 us01_U198 (.ZN( us01_n664 ) , .A1( us01_n726 ) , .A2( us01_n801 ) );
  OAI22_X1 us01_U199 (.ZN( us01_n708 ) , .A2( us01_n726 ) , .B2( us01_n727 ) , .A1( us01_n742 ) , .B1( us01_n811 ) );
  AOI222_X1 us01_U20 (.ZN( us01_n561 ) , .B1( us01_n828 ) , .C1( us01_n839 ) , .A2( us01_n841 ) , .A1( us01_n852 ) , .B2( us01_n861 ) , .C2( us01_n871 ) );
  NOR2_X1 us01_U200 (.ZN( us01_n650 ) , .A1( us01_n667 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U201 (.ZN( us01_n592 ) , .A2( us01_n695 ) , .A1( us01_n726 ) );
  NOR2_X1 us01_U202 (.A1( us01_n667 ) , .ZN( us01_n671 ) , .A2( us01_n742 ) );
  NOR2_X1 us01_U203 (.ZN( us01_n600 ) , .A1( us01_n667 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U204 (.A1( us01_n667 ) , .ZN( us01_n686 ) , .A2( us01_n814 ) );
  NOR2_X1 us01_U205 (.ZN( us01_n568 ) , .A1( us01_n726 ) , .A2( us01_n804 ) );
  NOR2_X1 us01_U206 (.A1( us01_n667 ) , .ZN( us01_n764 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U207 (.ZN( us01_n525 ) , .A1( us01_n667 ) , .A2( us01_n777 ) );
  NOR2_X1 us01_U208 (.ZN( us01_n652 ) , .A1( us01_n726 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U209 (.ZN( us01_n505 ) , .A1( us01_n810 ) , .A2( us01_n815 ) );
  NOR4_X1 us01_U21 (.ZN( us01_n471 ) , .A2( us01_n519 ) , .A4( us01_n592 ) , .A1( us01_n607 ) , .A3( us01_n627 ) );
  NOR2_X1 us01_U210 (.ZN( us01_n659 ) , .A1( us01_n727 ) , .A2( us01_n788 ) );
  NOR2_X1 us01_U211 (.ZN( us01_n544 ) , .A2( us01_n778 ) , .A1( us01_n812 ) );
  NOR2_X1 us01_U212 (.ZN( us01_n575 ) , .A2( us01_n697 ) , .A1( us01_n812 ) );
  NOR2_X1 us01_U213 (.ZN( us01_n507 ) , .A1( us01_n727 ) , .A2( us01_n777 ) );
  NOR2_X1 us01_U214 (.ZN( us01_n716 ) , .A2( us01_n722 ) , .A1( us01_n742 ) );
  INV_X1 us01_U215 (.A( us01_n748 ) , .ZN( us01_n840 ) );
  NOR2_X1 us01_U216 (.ZN( us01_n530 ) , .A2( us01_n747 ) , .A1( us01_n748 ) );
  NOR2_X1 us01_U217 (.ZN( us01_n660 ) , .A2( us01_n695 ) , .A1( us01_n727 ) );
  NOR2_X1 us01_U218 (.ZN( us01_n613 ) , .A1( us01_n783 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U219 (.ZN( us01_n627 ) , .A2( us01_n726 ) , .A1( us01_n783 ) );
  NOR4_X1 us01_U22 (.ZN( us01_n477 ) , .A1( us01_n518 ) , .A4( us01_n555 ) , .A3( us01_n580 ) , .A2( us01_n628 ) );
  NOR2_X1 us01_U220 (.ZN( us01_n609 ) , .A2( us01_n778 ) , .A1( us01_n804 ) );
  NOR2_X1 us01_U221 (.ZN( us01_n661 ) , .A1( us01_n727 ) , .A2( us01_n783 ) );
  NOR2_X1 us01_U222 (.ZN( us01_n626 ) , .A2( us01_n667 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U223 (.ZN( us01_n599 ) , .A2( us01_n778 ) , .A1( us01_n801 ) );
  INV_X1 us01_U224 (.A( us01_n745 ) , .ZN( us01_n832 ) );
  NOR2_X1 us01_U225 (.ZN( us01_n554 ) , .A1( us01_n760 ) , .A2( us01_n803 ) );
  NOR2_X1 us01_U226 (.ZN( us01_n529 ) , .A2( us01_n778 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U227 (.ZN( us01_n526 ) , .A2( us01_n722 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U228 (.A2( us01_n706 ) , .A1( us01_n748 ) , .ZN( us01_n769 ) );
  NOR2_X1 us01_U229 (.ZN( us01_n597 ) , .A2( us01_n789 ) , .A1( us01_n814 ) );
  NOR4_X1 us01_U23 (.ZN( us01_n454 ) , .A2( us01_n515 ) , .A1( us01_n541 ) , .A3( us01_n577 ) , .A4( us01_n613 ) );
  NOR2_X1 us01_U230 (.ZN( us01_n555 ) , .A1( us01_n790 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U231 (.ZN( us01_n542 ) , .A2( us01_n783 ) , .A1( us01_n790 ) );
  NOR2_X1 us01_U232 (.A2( us01_n695 ) , .ZN( us01_n714 ) , .A1( us01_n790 ) );
  NOR2_X1 us01_U233 (.ZN( us01_n665 ) , .A1( us01_n748 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U234 (.ZN( us01_n543 ) , .A1( us01_n747 ) , .A2( us01_n812 ) );
  NOR2_X1 us01_U235 (.ZN( us01_n553 ) , .A1( us01_n748 ) , .A2( us01_n789 ) );
  NOR2_X1 us01_U236 (.ZN( us01_n506 ) , .A2( us01_n778 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U237 (.ZN( us01_n541 ) , .A2( us01_n706 ) , .A1( us01_n783 ) );
  NOR2_X1 us01_U238 (.ZN( us01_n514 ) , .A1( us01_n706 ) , .A2( us01_n742 ) );
  NOR2_X1 us01_U239 (.ZN( us01_n662 ) , .A1( us01_n783 ) , .A2( us01_n789 ) );
  NOR4_X1 us01_U24 (.A4( us01_n530 ) , .A3( us01_n531 ) , .A2( us01_n532 ) , .ZN( us01_n533 ) , .A1( us01_n818 ) );
  NOR2_X1 us01_U240 (.ZN( us01_n556 ) , .A1( us01_n706 ) , .A2( us01_n814 ) );
  NOR2_X1 us01_U241 (.ZN( us01_n515 ) , .A1( us01_n706 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U242 (.ZN( us01_n612 ) , .A1( us01_n760 ) , .A2( us01_n810 ) );
  NOR2_X1 us01_U243 (.ZN( us01_n629 ) , .A1( us01_n722 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U244 (.A1( us01_n747 ) , .ZN( us01_n765 ) , .A2( us01_n801 ) );
  NOR2_X1 us01_U245 (.ZN( us01_n528 ) , .A2( us01_n742 ) , .A1( us01_n790 ) );
  INV_X1 us01_U246 (.A( us01_n804 ) , .ZN( us01_n839 ) );
  OAI22_X1 us01_U247 (.B1( us01_n438 ) , .ZN( us01_n442 ) , .A2( us01_n726 ) , .A1( us01_n742 ) , .B2( us01_n747 ) );
  NOR3_X1 us01_U248 (.ZN( us01_n438 ) , .A2( us01_n834 ) , .A3( us01_n835 ) , .A1( us01_n844 ) );
  INV_X1 us01_U249 (.A( us01_n726 ) , .ZN( us01_n850 ) );
  NOR4_X1 us01_U25 (.A4( us01_n539 ) , .A3( us01_n540 ) , .A2( us01_n541 ) , .ZN( us01_n548 ) , .A1( us01_n686 ) );
  NOR2_X1 us01_U250 (.ZN( us01_n519 ) , .A1( us01_n788 ) , .A2( us01_n810 ) );
  NOR2_X1 us01_U251 (.ZN( us01_n668 ) , .A1( us01_n788 ) , .A2( us01_n803 ) );
  AOI21_X1 us01_U252 (.ZN( us01_n550 ) , .B1( us01_n667 ) , .A( us01_n695 ) , .B2( us01_n803 ) );
  AOI21_X1 us01_U253 (.ZN( us01_n587 ) , .B2( us01_n697 ) , .B1( us01_n813 ) , .A( us01_n815 ) );
  NOR2_X1 us01_U254 (.ZN( us01_n504 ) , .A2( us01_n726 ) , .A1( us01_n760 ) );
  NOR2_X1 us01_U255 (.ZN( us01_n653 ) , .A1( us01_n788 ) , .A2( us01_n813 ) );
  INV_X1 us01_U256 (.A( us01_n801 ) , .ZN( us01_n841 ) );
  NOR2_X1 us01_U257 (.ZN( us01_n628 ) , .A1( us01_n745 ) , .A2( us01_n813 ) );
  NOR2_X1 us01_U258 (.ZN( us01_n545 ) , .A1( us01_n697 ) , .A2( us01_n742 ) );
  INV_X1 us01_U259 (.A( us01_n697 ) , .ZN( us01_n851 ) );
  NOR2_X1 us01_U26 (.ZN( us01_n678 ) , .A2( us01_n832 ) , .A1( us01_n837 ) );
  NOR2_X1 us01_U260 (.ZN( us01_n640 ) , .A2( us01_n786 ) , .A1( us01_n789 ) );
  AOI21_X1 us01_U261 (.ZN( us01_n648 ) , .A( us01_n777 ) , .B1( us01_n790 ) , .B2( us01_n803 ) );
  NOR2_X1 us01_U262 (.ZN( us01_n666 ) , .A2( us01_n706 ) , .A1( us01_n788 ) );
  NOR2_X1 us01_U263 (.A2( us01_n695 ) , .A1( us01_n778 ) , .ZN( us01_n818 ) );
  NOR2_X1 us01_U264 (.A1( us01_n695 ) , .ZN( us01_n768 ) , .A2( us01_n813 ) );
  AOI21_X1 us01_U265 (.ZN( us01_n624 ) , .B2( us01_n667 ) , .A( us01_n788 ) , .B1( us01_n789 ) );
  NOR2_X1 us01_U266 (.ZN( us01_n577 ) , .A2( us01_n706 ) , .A1( us01_n728 ) );
  INV_X1 us01_U267 (.A( us01_n761 ) , .ZN( us01_n864 ) );
  NOR2_X1 us01_U268 (.A2( us01_n706 ) , .A1( us01_n760 ) , .ZN( us01_n792 ) );
  NOR2_X1 us01_U269 (.ZN( us01_n607 ) , .A2( us01_n722 ) , .A1( us01_n815 ) );
  AOI222_X1 us01_U27 (.ZN( us01_n467 ) , .B1( us01_n830 ) , .A1( us01_n837 ) , .C1( us01_n840 ) , .C2( us01_n849 ) , .A2( us01_n853 ) , .B2( us01_n863 ) );
  NOR2_X1 us01_U270 (.ZN( us01_n531 ) , .A2( us01_n722 ) , .A1( us01_n728 ) );
  AOI21_X1 us01_U271 (.ZN( us01_n508 ) , .B2( us01_n667 ) , .A( us01_n728 ) , .B1( us01_n813 ) );
  AOI21_X1 us01_U272 (.ZN( us01_n537 ) , .B2( us01_n810 ) , .A( us01_n812 ) , .B1( us01_n813 ) );
  INV_X1 us01_U273 (.A( us01_n727 ) , .ZN( us01_n866 ) );
  NOR2_X1 us01_U274 (.ZN( us01_n540 ) , .A1( us01_n760 ) , .A2( us01_n789 ) );
  INV_X1 us01_U275 (.A( us01_n810 ) , .ZN( us01_n852 ) );
  AOI21_X1 us01_U276 (.B1( us01_n697 ) , .ZN( us01_n698 ) , .A( us01_n730 ) , .B2( us01_n761 ) );
  NOR2_X1 us01_U277 (.ZN( us01_n579 ) , .A1( us01_n667 ) , .A2( us01_n786 ) );
  AOI21_X1 us01_U278 (.ZN( us01_n589 ) , .B2( us01_n761 ) , .A( us01_n783 ) , .B1( us01_n810 ) );
  NOR2_X1 us01_U279 (.ZN( us01_n654 ) , .A1( us01_n745 ) , .A2( us01_n778 ) );
  NOR4_X1 us01_U28 (.A1( us01_n464 ) , .ZN( us01_n465 ) , .A4( us01_n540 ) , .A2( us01_n552 ) , .A3( us01_n612 ) );
  INV_X1 us01_U280 (.A( us01_n789 ) , .ZN( us01_n871 ) );
  AOI21_X1 us01_U281 (.B1( us01_n623 ) , .ZN( us01_n625 ) , .A( us01_n761 ) , .B2( us01_n812 ) );
  NOR2_X1 us01_U282 (.ZN( us01_n683 ) , .A1( us01_n727 ) , .A2( us01_n814 ) );
  AOI21_X1 us01_U283 (.A( us01_n813 ) , .B2( us01_n814 ) , .B1( us01_n815 ) , .ZN( us01_n816 ) );
  AOI21_X1 us01_U284 (.ZN( us01_n647 ) , .B1( us01_n727 ) , .B2( us01_n761 ) , .A( us01_n811 ) );
  AOI21_X1 us01_U285 (.A( us01_n810 ) , .B2( us01_n811 ) , .B1( us01_n812 ) , .ZN( us01_n817 ) );
  AOI21_X1 us01_U286 (.ZN( us01_n513 ) , .A( us01_n727 ) , .B1( us01_n748 ) , .B2( us01_n801 ) );
  AOI21_X1 us01_U287 (.ZN( us01_n497 ) , .B1( us01_n678 ) , .A( us01_n810 ) , .B2( us01_n814 ) );
  NOR2_X1 us01_U288 (.ZN( us01_n518 ) , .A2( us01_n706 ) , .A1( us01_n812 ) );
  AOI21_X1 us01_U289 (.ZN( us01_n475 ) , .A( us01_n667 ) , .B1( us01_n748 ) , .B2( us01_n804 ) );
  AOI221_X1 us01_U29 (.ZN( us01_n466 ) , .C2( us01_n712 ) , .B2( us01_n829 ) , .C1( us01_n843 ) , .B1( us01_n858 ) , .A( us01_n862 ) );
  NOR2_X1 us01_U290 (.ZN( us01_n566 ) , .A1( us01_n727 ) , .A2( us01_n760 ) );
  NOR2_X1 us01_U291 (.ZN( us01_n580 ) , .A1( us01_n742 ) , .A2( us01_n813 ) );
  AOI21_X1 us01_U292 (.ZN( us01_n591 ) , .B1( us01_n748 ) , .A( us01_n790 ) , .B2( us01_n811 ) );
  NOR2_X1 us01_U293 (.ZN( us01_n564 ) , .A2( us01_n695 ) , .A1( us01_n761 ) );
  AOI21_X1 us01_U294 (.ZN( us01_n512 ) , .A( us01_n777 ) , .B2( us01_n790 ) , .B1( us01_n810 ) );
  NAND2_X2 us01_U295 (.A2( us01_n462 ) , .A1( us01_n463 ) , .ZN( us01_n810 ) );
  AOI21_X1 us01_U296 (.ZN( us01_n637 ) , .B2( us01_n747 ) , .A( us01_n786 ) , .B1( us01_n810 ) );
  NOR2_X1 us01_U297 (.ZN( us01_n557 ) , .A2( us01_n789 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U298 (.A2( us01_n811 ) , .A1( us01_n813 ) , .ZN( us01_n819 ) );
  NOR2_X1 us01_U299 (.ZN( us01_n527 ) , .A1( us01_n706 ) , .A2( us01_n777 ) );
  NAND2_X2 us01_U3 (.A1( us01_n447 ) , .A2( us01_n462 ) , .ZN( us01_n722 ) );
  NOR4_X1 us01_U30 (.A4( us01_n512 ) , .A3( us01_n513 ) , .A2( us01_n514 ) , .A1( us01_n515 ) , .ZN( us01_n522 ) );
  NOR2_X1 us01_U300 (.ZN( us01_n517 ) , .A2( us01_n697 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U301 (.ZN( us01_n681 ) , .A2( us01_n697 ) , .A1( us01_n801 ) );
  NOR2_X1 us01_U302 (.ZN( us01_n576 ) , .A1( us01_n706 ) , .A2( us01_n811 ) );
  INV_X1 us01_U303 (.A( us01_n813 ) , .ZN( us01_n853 ) );
  INV_X1 us01_U304 (.A( us01_n811 ) , .ZN( us01_n834 ) );
  AOI21_X1 us01_U305 (.ZN( us01_n448 ) , .B2( us01_n790 ) , .A( us01_n801 ) , .B1( us01_n813 ) );
  AOI21_X1 us01_U306 (.ZN( us01_n538 ) , .A( us01_n761 ) , .B2( us01_n777 ) , .B1( us01_n815 ) );
  AOI21_X1 us01_U307 (.ZN( us01_n496 ) , .A( us01_n722 ) , .B2( us01_n760 ) , .B1( us01_n812 ) );
  AOI21_X1 us01_U308 (.ZN( us01_n687 ) , .B2( us01_n747 ) , .B1( us01_n761 ) , .A( us01_n804 ) );
  AOI21_X1 us01_U309 (.B1( us01_n684 ) , .ZN( us01_n685 ) , .A( us01_n726 ) , .B2( us01_n759 ) );
  AOI222_X1 us01_U31 (.ZN( us01_n523 ) , .A1( us01_n832 ) , .B2( us01_n835 ) , .C1( us01_n842 ) , .C2( us01_n848 ) , .A2( us01_n850 ) , .B1( us01_n864 ) );
  NOR2_X1 us01_U310 (.ZN( us01_n581 ) , .A1( us01_n790 ) , .A2( us01_n815 ) );
  NOR2_X1 us01_U311 (.ZN( us01_n532 ) , .A1( us01_n722 ) , .A2( us01_n786 ) );
  NOR2_X1 us01_U312 (.ZN( us01_n630 ) , .A2( us01_n695 ) , .A1( us01_n722 ) );
  AOI21_X1 us01_U313 (.A( us01_n788 ) , .B2( us01_n789 ) , .B1( us01_n790 ) , .ZN( us01_n791 ) );
  AOI21_X1 us01_U314 (.A( us01_n731 ) , .ZN( us01_n732 ) , .B2( us01_n778 ) , .B1( us01_n790 ) );
  NOR2_X1 us01_U315 (.ZN( us01_n565 ) , .A1( us01_n745 ) , .A2( us01_n803 ) );
  AOI21_X1 us01_U316 (.ZN( us01_n567 ) , .B1( us01_n748 ) , .B2( us01_n760 ) , .A( us01_n778 ) );
  AOI21_X1 us01_U317 (.ZN( us01_n638 ) , .B2( us01_n745 ) , .A( us01_n790 ) , .B1( us01_n801 ) );
  AOI21_X1 us01_U318 (.ZN( us01_n562 ) , .B1( us01_n722 ) , .A( us01_n777 ) , .B2( us01_n789 ) );
  AOI21_X1 us01_U319 (.ZN( us01_n569 ) , .B2( us01_n695 ) , .B1( us01_n804 ) , .A( us01_n810 ) );
  NOR4_X1 us01_U32 (.A3( us01_n519 ) , .A1( us01_n520 ) , .ZN( us01_n521 ) , .A2( us01_n671 ) , .A4( us01_n767 ) );
  NOR2_X1 us01_U320 (.ZN( us01_n663 ) , .A1( us01_n778 ) , .A2( us01_n811 ) );
  NOR2_X1 us01_U321 (.ZN( us01_n578 ) , .A2( us01_n695 ) , .A1( us01_n789 ) );
  NOR2_X1 us01_U322 (.ZN( us01_n682 ) , .A1( us01_n789 ) , .A2( us01_n811 ) );
  NAND2_X2 us01_U323 (.A1( us01_n450 ) , .A2( us01_n463 ) , .ZN( us01_n667 ) );
  NAND2_X1 us01_U324 (.ZN( us01_n751 ) , .A1( us01_n761 ) , .A2( us01_n803 ) );
  NOR2_X1 us01_U325 (.ZN( us01_n709 ) , .A1( us01_n760 ) , .A2( us01_n761 ) );
  AOI21_X1 us01_U326 (.ZN( us01_n476 ) , .B2( us01_n695 ) , .A( us01_n747 ) , .B1( us01_n777 ) );
  NOR2_X1 us01_U327 (.ZN( us01_n680 ) , .A2( us01_n706 ) , .A1( us01_n815 ) );
  INV_X1 us01_U328 (.A( us01_n778 ) , .ZN( us01_n848 ) );
  OAI21_X1 us01_U329 (.A( us01_n729 ) , .B1( us01_n730 ) , .ZN( us01_n734 ) , .B2( us01_n803 ) );
  AOI221_X1 us01_U33 (.A( us01_n779 ) , .ZN( us01_n796 ) , .C2( us01_n835 ) , .B2( us01_n836 ) , .B1( us01_n863 ) , .C1( us01_n864 ) );
  OAI21_X1 us01_U330 (.ZN( us01_n729 ) , .A( us01_n831 ) , .B2( us01_n850 ) , .B1( us01_n871 ) );
  AOI21_X1 us01_U331 (.ZN( us01_n639 ) , .B1( us01_n678 ) , .A( us01_n789 ) , .B2( us01_n815 ) );
  AOI21_X1 us01_U332 (.ZN( us01_n440 ) , .A( us01_n697 ) , .B1( us01_n731 ) , .B2( us01_n748 ) );
  NAND2_X1 us01_U333 (.A1( us01_n697 ) , .A2( us01_n727 ) , .ZN( us01_n780 ) );
  NOR2_X1 us01_U334 (.ZN( us01_n468 ) , .A2( us01_n777 ) , .A1( us01_n813 ) );
  NOR2_X1 us01_U335 (.ZN( us01_n516 ) , .A1( us01_n706 ) , .A2( us01_n786 ) );
  NAND2_X2 us01_U336 (.A2( us01_n447 ) , .A1( us01_n450 ) , .ZN( us01_n761 ) );
  OAI21_X1 us01_U337 (.A( us01_n696 ) , .ZN( us01_n700 ) , .B2( us01_n748 ) , .B1( us01_n802 ) );
  OAI21_X1 us01_U338 (.ZN( us01_n696 ) , .B2( us01_n831 ) , .B1( us01_n836 ) , .A( us01_n858 ) );
  NOR2_X1 us01_U339 (.ZN( us01_n524 ) , .A1( us01_n722 ) , .A2( us01_n748 ) );
  NOR4_X1 us01_U34 (.A4( us01_n791 ) , .A3( us01_n792 ) , .A2( us01_n793 ) , .A1( us01_n794 ) , .ZN( us01_n795 ) );
  AOI21_X1 us01_U340 (.ZN( us01_n441 ) , .B1( us01_n787 ) , .B2( us01_n789 ) , .A( us01_n812 ) );
  AOI21_X1 us01_U341 (.ZN( us01_n495 ) , .A( us01_n777 ) , .B2( us01_n789 ) , .B1( us01_n802 ) );
  NAND2_X1 us01_U342 (.ZN( us01_n712 ) , .A1( us01_n726 ) , .A2( us01_n778 ) );
  NOR2_X1 us01_U343 (.ZN( us01_n482 ) , .A1( us01_n786 ) , .A2( us01_n803 ) );
  NAND2_X1 us01_U344 (.A2( us01_n760 ) , .A1( us01_n804 ) , .ZN( us01_n808 ) );
  OAI21_X1 us01_U345 (.A( us01_n785 ) , .B2( us01_n786 ) , .B1( us01_n787 ) , .ZN( us01_n793 ) );
  OAI21_X1 us01_U346 (.ZN( us01_n785 ) , .A( us01_n837 ) , .B1( us01_n861 ) , .B2( us01_n871 ) );
  INV_X1 us01_U347 (.A( us01_n783 ) , .ZN( us01_n844 ) );
  NOR2_X1 us01_U348 (.ZN( us01_n710 ) , .A2( us01_n722 ) , .A1( us01_n788 ) );
  NAND2_X1 us01_U349 (.ZN( us01_n669 ) , .A1( us01_n804 ) , .A2( us01_n814 ) );
  NOR4_X1 us01_U35 (.A4( us01_n774 ) , .A3( us01_n775 ) , .A1( us01_n776 ) , .ZN( us01_n797 ) , .A2( us01_n799 ) );
  NAND2_X2 us01_U350 (.A2( us01_n446 ) , .A1( us01_n450 ) , .ZN( us01_n727 ) );
  INV_X1 us01_U351 (.A( us01_n722 ) , .ZN( us01_n854 ) );
  NAND2_X2 us01_U352 (.A1( us01_n445 ) , .A2( us01_n463 ) , .ZN( us01_n747 ) );
  INV_X1 us01_U353 (.A( us01_n815 ) , .ZN( us01_n842 ) );
  AND2_X1 us01_U354 (.ZN( us01_n730 ) , .A1( us01_n777 ) , .A2( us01_n783 ) );
  NAND2_X1 us01_U355 (.A1( us01_n445 ) , .A2( us01_n447 ) , .ZN( us01_n803 ) );
  NAND2_X1 us01_U356 (.A1( us01_n449 ) , .A2( us01_n452 ) , .ZN( us01_n812 ) );
  NAND2_X1 us01_U357 (.A1( us01_n453 ) , .A2( us01_n469 ) , .ZN( us01_n801 ) );
  NAND2_X1 us01_U358 (.A1( us01_n453 ) , .A2( us01_n460 ) , .ZN( us01_n748 ) );
  NAND2_X2 us01_U359 (.A2( us01_n446 ) , .A1( us01_n458 ) , .ZN( us01_n726 ) );
  NOR2_X1 us01_U36 (.ZN( us01_n802 ) , .A1( us01_n852 ) , .A2( us01_n859 ) );
  NAND2_X1 us01_U360 (.A2( us01_n451 ) , .A1( us01_n453 ) , .ZN( us01_n804 ) );
  NAND2_X1 us01_U361 (.A1( us01_n449 ) , .A2( us01_n469 ) , .ZN( us01_n814 ) );
  NAND2_X1 us01_U362 (.A1( us01_n452 ) , .A2( us01_n459 ) , .ZN( us01_n811 ) );
  NAND2_X1 us01_U363 (.A1( us01_n451 ) , .A2( us01_n459 ) , .ZN( us01_n742 ) );
  NAND2_X1 us01_U364 (.A1( us01_n451 ) , .A2( us01_n470 ) , .ZN( us01_n783 ) );
  NAND2_X1 us01_U365 (.A2( us01_n452 ) , .A1( us01_n470 ) , .ZN( us01_n777 ) );
  NAND2_X1 us01_U366 (.A2( us01_n459 ) , .A1( us01_n460 ) , .ZN( us01_n745 ) );
  NAND2_X2 us01_U367 (.A2( us01_n446 ) , .A1( us01_n462 ) , .ZN( us01_n813 ) );
  NAND2_X1 us01_U368 (.A1( us01_n460 ) , .A2( us01_n470 ) , .ZN( us01_n786 ) );
  NOR2_X1 us01_U369 (.ZN( us01_n451 ) , .A1( us01_n824 ) , .A2( us01_n825 ) );
  NAND4_X1 us01_U37 (.ZN( sa01_sr_2 ) , .A4( us01_n641 ) , .A3( us01_n642 ) , .A2( us01_n643 ) , .A1( us01_n644 ) );
  NOR2_X1 us01_U370 (.ZN( us01_n449 ) , .A1( us01_n826 ) , .A2( us01_n827 ) );
  NAND2_X1 us01_U371 (.A1( us01_n449 ) , .A2( us01_n460 ) , .ZN( us01_n788 ) );
  NAND2_X2 us01_U372 (.A1( us01_n447 ) , .A2( us01_n458 ) , .ZN( us01_n790 ) );
  NAND2_X2 us01_U373 (.A2( us01_n439 ) , .A1( us01_n450 ) , .ZN( us01_n789 ) );
  NAND2_X1 us01_U374 (.A2( us01_n452 ) , .A1( us01_n453 ) , .ZN( us01_n728 ) );
  NAND2_X2 us01_U375 (.A2( us01_n469 ) , .A1( us01_n470 ) , .ZN( us01_n815 ) );
  NAND2_X1 us01_U376 (.A1( us01_n445 ) , .A2( us01_n446 ) , .ZN( us01_n784 ) );
  NAND2_X2 us01_U377 (.A2( us01_n439 ) , .A1( us01_n445 ) , .ZN( us01_n782 ) );
  NOR2_X1 us01_U378 (.A2( sa01_7 ) , .ZN( us01_n458 ) , .A1( us01_n847 ) );
  NOR2_X1 us01_U379 (.A2( sa01_2 ) , .A1( sa01_3 ) , .ZN( us01_n470 ) );
  AOI222_X1 us01_U38 (.B2( us01_n636 ) , .ZN( us01_n642 ) , .B1( us01_n839 ) , .A1( us01_n840 ) , .C2( us01_n844 ) , .C1( us01_n861 ) , .A2( us01_n863 ) );
  NOR2_X1 us01_U380 (.A2( sa01_1 ) , .ZN( us01_n469 ) , .A1( us01_n824 ) );
  NOR2_X1 us01_U381 (.A2( sa01_0 ) , .ZN( us01_n452 ) , .A1( us01_n825 ) );
  NOR2_X1 us01_U382 (.A2( sa01_0 ) , .A1( sa01_1 ) , .ZN( us01_n460 ) );
  NAND2_X2 us01_U383 (.A1( us01_n439 ) , .A2( us01_n458 ) , .ZN( us01_n697 ) );
  NOR2_X1 us01_U384 (.A2( sa01_3 ) , .ZN( us01_n453 ) , .A1( us01_n826 ) );
  NOR2_X1 us01_U385 (.A2( sa01_2 ) , .ZN( us01_n459 ) , .A1( us01_n827 ) );
  INV_X1 us01_U386 (.A( sa01_3 ) , .ZN( us01_n827 ) );
  INV_X1 us01_U387 (.A( sa01_1 ) , .ZN( us01_n825 ) );
  INV_X1 us01_U388 (.A( sa01_0 ) , .ZN( us01_n824 ) );
  INV_X1 us01_U389 (.A( sa01_2 ) , .ZN( us01_n826 ) );
  NOR4_X1 us01_U39 (.A4( us01_n637 ) , .A3( us01_n638 ) , .A2( us01_n639 ) , .A1( us01_n640 ) , .ZN( us01_n641 ) );
  INV_X1 us01_U390 (.A( sa01_5 ) , .ZN( us01_n846 ) );
  NAND2_X1 us01_U391 (.A1( us01_n727 ) , .A2( us01_n782 ) , .ZN( us01_n809 ) );
  OAI22_X1 us01_U392 (.ZN( us01_n586 ) , .A2( us01_n745 ) , .B2( us01_n760 ) , .A1( us01_n761 ) , .B1( us01_n782 ) );
  AOI21_X1 us01_U393 (.ZN( us01_n590 ) , .B1( us01_n726 ) , .B2( us01_n782 ) , .A( us01_n788 ) );
  AOI21_X1 us01_U394 (.ZN( us01_n646 ) , .A( us01_n760 ) , .B2( us01_n782 ) , .B1( us01_n790 ) );
  AOI21_X1 us01_U395 (.ZN( us01_n621 ) , .B1( us01_n697 ) , .A( us01_n777 ) , .B2( us01_n782 ) );
  OAI22_X1 us01_U396 (.ZN( us01_n679 ) , .A1( us01_n697 ) , .A2( us01_n728 ) , .B2( us01_n782 ) , .B1( us01_n815 ) );
  OAI21_X1 us01_U397 (.A( us01_n611 ) , .ZN( us01_n614 ) , .B1( us01_n623 ) , .B2( us01_n782 ) );
  NOR2_X1 us01_U398 (.ZN( us01_n608 ) , .A1( us01_n782 ) , .A2( us01_n814 ) );
  INV_X2 us01_U399 (.A( us01_n747 ) , .ZN( us01_n861 ) );
  NAND2_X2 us01_U4 (.A1( us01_n439 ) , .A2( us01_n462 ) , .ZN( us01_n706 ) );
  NOR3_X1 us01_U40 (.A2( us01_n605 ) , .A1( us01_n606 ) , .ZN( us01_n644 ) , .A3( us01_n720 ) );
  OAI222_X1 us01_U400 (.A2( us01_n667 ) , .ZN( us01_n672 ) , .B1( us01_n745 ) , .B2( us01_n782 ) , .C2( us01_n786 ) , .C1( us01_n813 ) , .A1( us01_n815 ) );
  NOR2_X1 us01_U401 (.ZN( us01_n649 ) , .A1( us01_n782 ) , .A2( us01_n786 ) );
  NOR2_X1 us01_U402 (.ZN( us01_n598 ) , .A2( us01_n695 ) , .A1( us01_n782 ) );
  NOR2_X1 us01_U403 (.ZN( us01_n551 ) , .A2( us01_n742 ) , .A1( us01_n782 ) );
  INV_X1 us01_U404 (.A( us01_n782 ) , .ZN( us01_n859 ) );
  NAND2_X1 us01_U405 (.A2( us01_n459 ) , .A1( us01_n469 ) , .ZN( us01_n695 ) );
  INV_X1 us01_U406 (.A( sa01_7 ) , .ZN( us01_n856 ) );
  OAI221_X1 us01_U407 (.A( us01_n781 ) , .C2( us01_n782 ) , .B2( us01_n783 ) , .B1( us01_n784 ) , .ZN( us01_n794 ) , .C1( us01_n811 ) );
  AOI21_X1 us01_U408 (.ZN( us01_n498 ) , .A( us01_n695 ) , .B1( us01_n706 ) , .B2( us01_n784 ) );
  OAI221_X1 us01_U409 (.A( us01_n694 ) , .ZN( us01_n701 ) , .C2( us01_n782 ) , .C1( us01_n783 ) , .B1( us01_n784 ) , .B2( us01_n804 ) );
  NAND4_X1 us01_U41 (.ZN( sa01_sr_7 ) , .A4( us01_n820 ) , .A3( us01_n821 ) , .A2( us01_n822 ) , .A1( us01_n823 ) );
  OAI22_X1 us01_U410 (.ZN( us01_n588 ) , .B1( us01_n728 ) , .B2( us01_n747 ) , .A2( us01_n784 ) , .A1( us01_n801 ) );
  AOI222_X1 us01_U411 (.ZN( us01_n511 ) , .C1( us01_n830 ) , .B2( us01_n835 ) , .A2( us01_n841 ) , .C2( us01_n860 ) , .B1( us01_n861 ) , .A1( us01_n864 ) );
  AOI222_X1 us01_U412 (.ZN( us01_n603 ) , .B2( us01_n669 ) , .B1( us01_n751 ) , .C2( us01_n829 ) , .A1( us01_n831 ) , .A2( us01_n860 ) , .C1( us01_n861 ) );
  AOI221_X1 us01_U413 (.A( us01_n481 ) , .ZN( us01_n486 ) , .B1( us01_n829 ) , .C2( us01_n842 ) , .C1( us01_n850 ) , .B2( us01_n860 ) );
  NAND2_X1 us01_U414 (.A2( us01_n747 ) , .A1( us01_n784 ) , .ZN( us01_n807 ) );
  NOR2_X1 us01_U415 (.ZN( us01_n610 ) , .A1( us01_n777 ) , .A2( us01_n784 ) );
  NOR2_X1 us01_U416 (.ZN( us01_n715 ) , .A2( us01_n742 ) , .A1( us01_n784 ) );
  OAI222_X1 us01_U417 (.ZN( us01_n615 ) , .B1( us01_n695 ) , .C1( us01_n722 ) , .C2( us01_n745 ) , .B2( us01_n784 ) , .A2( us01_n790 ) , .A1( us01_n814 ) );
  NOR2_X1 us01_U418 (.ZN( us01_n651 ) , .A1( us01_n760 ) , .A2( us01_n784 ) );
  NOR2_X1 us01_U419 (.ZN( us01_n552 ) , .A1( us01_n784 ) , .A2( us01_n811 ) );
  AOI222_X1 us01_U42 (.C2( us01_n807 ) , .B2( us01_n808 ) , .A2( us01_n809 ) , .ZN( us01_n821 ) , .C1( us01_n830 ) , .A1( us01_n837 ) , .B1( us01_n851 ) );
  NOR2_X1 us01_U420 (.ZN( us01_n787 ) , .A2( us01_n860 ) , .A1( us01_n866 ) );
  NOR2_X1 us01_U421 (.ZN( us01_n699 ) , .A2( us01_n784 ) , .A1( us01_n815 ) );
  NOR2_X1 us01_U422 (.A1( us01_n728 ) , .ZN( us01_n763 ) , .A2( us01_n784 ) );
  INV_X1 us01_U423 (.A( us01_n784 ) , .ZN( us01_n860 ) );
  NOR2_X1 us01_U424 (.A2( sa01_4 ) , .ZN( us01_n447 ) , .A1( us01_n846 ) );
  NOR2_X1 us01_U425 (.ZN( us01_n463 ) , .A2( us01_n845 ) , .A1( us01_n846 ) );
  NOR2_X1 us01_U426 (.A2( sa01_5 ) , .ZN( us01_n446 ) , .A1( us01_n845 ) );
  NOR2_X1 us01_U427 (.A2( sa01_4 ) , .A1( sa01_5 ) , .ZN( us01_n439 ) );
  INV_X1 us01_U428 (.A( sa01_6 ) , .ZN( us01_n847 ) );
  NOR2_X1 us01_U429 (.ZN( us01_n445 ) , .A2( us01_n847 ) , .A1( us01_n856 ) );
  NOR4_X1 us01_U43 (.A4( us01_n816 ) , .A3( us01_n817 ) , .A2( us01_n818 ) , .A1( us01_n819 ) , .ZN( us01_n820 ) );
  NOR2_X1 us01_U430 (.A2( sa01_6 ) , .ZN( us01_n450 ) , .A1( us01_n856 ) );
  NOR2_X1 us01_U431 (.A2( sa01_6 ) , .A1( sa01_7 ) , .ZN( us01_n462 ) );
  AOI221_X1 us01_U432 (.A( us01_n574 ) , .ZN( us01_n585 ) , .B2( us01_n829 ) , .C2( us01_n841 ) , .B1( us01_n852 ) , .C1( us01_n859 ) );
  AOI21_X1 us01_U433 (.ZN( us01_n574 ) , .B2( us01_n722 ) , .B1( us01_n746 ) , .A( us01_n783 ) );
  INV_X1 us01_U434 (.A( sa01_4 ) , .ZN( us01_n845 ) );
  AOI211_X1 us01_U435 (.A( us01_n635 ) , .ZN( us01_n643 ) , .B( us01_n741 ) , .C2( us01_n837 ) , .C1( us01_n852 ) );
  NAND4_X1 us01_U436 (.A4( us01_n631 ) , .A3( us01_n632 ) , .A2( us01_n633 ) , .A1( us01_n634 ) , .ZN( us01_n741 ) );
  NAND3_X1 us01_U437 (.ZN( sa01_sr_6 ) , .A3( us01_n795 ) , .A2( us01_n796 ) , .A1( us01_n797 ) );
  NAND3_X1 us01_U438 (.ZN( sa01_sr_5 ) , .A3( us01_n756 ) , .A2( us01_n757 ) , .A1( us01_n758 ) );
  NAND3_X1 us01_U439 (.ZN( sa01_sr_4 ) , .A3( us01_n736 ) , .A2( us01_n737 ) , .A1( us01_n738 ) );
  AOI211_X1 us01_U44 (.B( us01_n805 ) , .A( us01_n806 ) , .ZN( us01_n822 ) , .C1( us01_n840 ) , .C2( us01_n848 ) );
  NAND3_X1 us01_U440 (.A3( us01_n673 ) , .A2( us01_n674 ) , .A1( us01_n675 ) , .ZN( us01_n805 ) );
  NAND3_X1 us01_U441 (.ZN( us01_n636 ) , .A3( us01_n706 ) , .A2( us01_n722 ) , .A1( us01_n790 ) );
  NAND3_X1 us01_U442 (.A3( us01_n616 ) , .A2( us01_n617 ) , .A1( us01_n618 ) , .ZN( us01_n723 ) );
  NAND3_X1 us01_U443 (.A3( us01_n583 ) , .A2( us01_n584 ) , .A1( us01_n585 ) , .ZN( us01_n619 ) );
  NAND3_X1 us01_U444 (.ZN( us01_n563 ) , .A3( us01_n678 ) , .A2( us01_n748 ) , .A1( us01_n783 ) );
  NAND3_X1 us01_U445 (.A3( us01_n521 ) , .A2( us01_n522 ) , .A1( us01_n523 ) , .ZN( us01_n740 ) );
  NAND3_X1 us01_U446 (.A3( us01_n510 ) , .A1( us01_n511 ) , .ZN( us01_n606 ) , .A2( us01_n869 ) );
  NAND3_X1 us01_U447 (.A3( us01_n465 ) , .A2( us01_n466 ) , .A1( us01_n467 ) , .ZN( us01_n775 ) );
  NAND4_X1 us01_U45 (.ZN( sa01_sr_0 ) , .A4( us01_n499 ) , .A3( us01_n500 ) , .A2( us01_n501 ) , .A1( us01_n502 ) );
  NOR4_X1 us01_U46 (.A4( us01_n496 ) , .A3( us01_n497 ) , .A2( us01_n498 ) , .ZN( us01_n499 ) , .A1( us01_n525 ) );
  AOI221_X1 us01_U47 (.A( us01_n495 ) , .ZN( us01_n500 ) , .B2( us01_n841 ) , .C1( us01_n844 ) , .C2( us01_n858 ) , .B1( us01_n860 ) );
  AOI211_X1 us01_U48 (.A( us01_n494 ) , .ZN( us01_n501 ) , .B( us01_n800 ) , .C2( us01_n837 ) , .C1( us01_n849 ) );
  NOR2_X1 us01_U49 (.ZN( us01_n746 ) , .A1( us01_n859 ) , .A2( us01_n860 ) );
  NAND2_X2 us01_U5 (.A2( us01_n458 ) , .A1( us01_n463 ) , .ZN( us01_n778 ) );
  NAND4_X1 us01_U50 (.ZN( sa01_sr_1 ) , .A4( us01_n593 ) , .A3( us01_n594 ) , .A2( us01_n595 ) , .A1( us01_n596 ) );
  AOI211_X1 us01_U51 (.B( us01_n587 ) , .A( us01_n588 ) , .ZN( us01_n594 ) , .C2( us01_n809 ) , .C1( us01_n831 ) );
  NOR4_X1 us01_U52 (.A4( us01_n589 ) , .A3( us01_n590 ) , .A2( us01_n591 ) , .A1( us01_n592 ) , .ZN( us01_n593 ) );
  AOI211_X1 us01_U53 (.A( us01_n586 ) , .ZN( us01_n595 ) , .B( us01_n619 ) , .C1( us01_n843 ) , .C2( us01_n853 ) );
  NOR2_X1 us01_U54 (.ZN( us01_n623 ) , .A2( us01_n834 ) , .A1( us01_n837 ) );
  NAND4_X1 us01_U55 (.A4( us01_n601 ) , .A3( us01_n602 ) , .A2( us01_n603 ) , .A1( us01_n604 ) , .ZN( us01_n720 ) );
  NOR3_X1 us01_U56 (.A1( us01_n597 ) , .ZN( us01_n602 ) , .A3( us01_n661 ) , .A2( us01_n768 ) );
  NOR4_X1 us01_U57 (.A3( us01_n598 ) , .A2( us01_n599 ) , .A1( us01_n600 ) , .ZN( us01_n601 ) , .A4( us01_n653 ) );
  AOI222_X1 us01_U58 (.ZN( us01_n604 ) , .A1( us01_n828 ) , .C2( us01_n835 ) , .B1( us01_n840 ) , .A2( us01_n854 ) , .B2( us01_n859 ) , .C1( us01_n866 ) );
  NOR4_X1 us01_U59 (.A4( us01_n575 ) , .A3( us01_n576 ) , .A2( us01_n577 ) , .ZN( us01_n584 ) , .A1( us01_n681 ) );
  INV_X1 us01_U6 (.A( us01_n667 ) , .ZN( us01_n863 ) );
  NOR4_X1 us01_U60 (.A1( us01_n582 ) , .ZN( us01_n583 ) , .A3( us01_n650 ) , .A2( us01_n660 ) , .A4( us01_n765 ) );
  NAND4_X1 us01_U61 (.A4( us01_n483 ) , .A3( us01_n484 ) , .A2( us01_n485 ) , .A1( us01_n486 ) , .ZN( us01_n776 ) );
  NOR4_X1 us01_U62 (.A4( us01_n482 ) , .ZN( us01_n485 ) , .A1( us01_n564 ) , .A2( us01_n579 ) , .A3( us01_n600 ) );
  NOR4_X1 us01_U63 (.ZN( us01_n483 ) , .A2( us01_n531 ) , .A1( us01_n556 ) , .A3( us01_n629 ) , .A4( us01_n716 ) );
  NOR4_X1 us01_U64 (.ZN( us01_n484 ) , .A1( us01_n505 ) , .A2( us01_n517 ) , .A4( us01_n544 ) , .A3( us01_n609 ) );
  NOR4_X1 us01_U65 (.A4( us01_n627 ) , .A3( us01_n628 ) , .A2( us01_n629 ) , .A1( us01_n630 ) , .ZN( us01_n631 ) );
  AOI211_X1 us01_U66 (.B( us01_n621 ) , .A( us01_n622 ) , .ZN( us01_n633 ) , .C2( us01_n834 ) , .C1( us01_n861 ) );
  NOR4_X1 us01_U67 (.A4( us01_n624 ) , .A3( us01_n625 ) , .A2( us01_n626 ) , .ZN( us01_n632 ) , .A1( us01_n662 ) );
  NAND4_X1 us01_U68 (.A4( us01_n655 ) , .A3( us01_n656 ) , .A2( us01_n657 ) , .A1( us01_n658 ) , .ZN( us01_n798 ) );
  NOR3_X1 us01_U69 (.A3( us01_n649 ) , .A2( us01_n650 ) , .A1( us01_n651 ) , .ZN( us01_n656 ) );
  NOR3_X1 us01_U7 (.ZN( us01_n596 ) , .A1( us01_n606 ) , .A3( us01_n721 ) , .A2( us01_n740 ) );
  NOR3_X1 us01_U70 (.A3( us01_n652 ) , .A2( us01_n653 ) , .A1( us01_n654 ) , .ZN( us01_n655 ) );
  NOR3_X1 us01_U71 (.A3( us01_n646 ) , .A2( us01_n647 ) , .A1( us01_n648 ) , .ZN( us01_n657 ) );
  NAND4_X1 us01_U72 (.A4( us01_n558 ) , .A3( us01_n559 ) , .A2( us01_n560 ) , .A1( us01_n561 ) , .ZN( us01_n605 ) );
  NOR4_X1 us01_U73 (.ZN( us01_n559 ) , .A1( us01_n651 ) , .A3( us01_n659 ) , .A4( us01_n683 ) , .A2( us01_n766 ) );
  NOR4_X1 us01_U74 (.A4( us01_n550 ) , .A3( us01_n551 ) , .A2( us01_n552 ) , .A1( us01_n553 ) , .ZN( us01_n560 ) );
  NOR4_X1 us01_U75 (.A4( us01_n554 ) , .A3( us01_n555 ) , .A2( us01_n556 ) , .A1( us01_n557 ) , .ZN( us01_n558 ) );
  NAND4_X1 us01_U76 (.A4( us01_n770 ) , .A3( us01_n771 ) , .A2( us01_n772 ) , .A1( us01_n773 ) , .ZN( us01_n799 ) );
  NOR3_X1 us01_U77 (.A3( us01_n763 ) , .A2( us01_n764 ) , .A1( us01_n765 ) , .ZN( us01_n771 ) );
  NOR4_X1 us01_U78 (.A4( us01_n766 ) , .A3( us01_n767 ) , .A2( us01_n768 ) , .A1( us01_n769 ) , .ZN( us01_n770 ) );
  AOI222_X1 us01_U79 (.ZN( us01_n773 ) , .A1( us01_n828 ) , .C1( us01_n832 ) , .B2( us01_n839 ) , .A2( us01_n848 ) , .B1( us01_n859 ) , .C2( us01_n871 ) );
  NOR3_X1 us01_U8 (.A3( us01_n798 ) , .A2( us01_n799 ) , .A1( us01_n800 ) , .ZN( us01_n823 ) );
  NOR4_X1 us01_U80 (.A4( us01_n507 ) , .A2( us01_n508 ) , .A1( us01_n509 ) , .ZN( us01_n510 ) , .A3( us01_n668 ) );
  INV_X1 us01_U81 (.A( us01_n503 ) , .ZN( us01_n869 ) );
  NOR4_X1 us01_U82 (.A4( us01_n663 ) , .A3( us01_n664 ) , .A2( us01_n665 ) , .A1( us01_n666 ) , .ZN( us01_n674 ) );
  NOR4_X1 us01_U83 (.A4( us01_n659 ) , .A3( us01_n660 ) , .A2( us01_n661 ) , .A1( us01_n662 ) , .ZN( us01_n675 ) );
  NOR4_X1 us01_U84 (.A3( us01_n671 ) , .A1( us01_n672 ) , .ZN( us01_n673 ) , .A4( us01_n713 ) , .A2( us01_n857 ) );
  NOR2_X1 us01_U85 (.ZN( us01_n759 ) , .A1( us01_n831 ) , .A2( us01_n832 ) );
  NAND4_X1 us01_U86 (.A4( us01_n454 ) , .A3( us01_n455 ) , .A2( us01_n456 ) , .A1( us01_n457 ) , .ZN( us01_n677 ) );
  NOR3_X1 us01_U87 (.ZN( us01_n455 ) , .A3( us01_n528 ) , .A1( us01_n553 ) , .A2( us01_n568 ) );
  AOI221_X1 us01_U88 (.A( us01_n448 ) , .ZN( us01_n457 ) , .C2( us01_n751 ) , .B1( us01_n830 ) , .C1( us01_n840 ) , .B2( us01_n859 ) );
  NOR4_X1 us01_U89 (.ZN( us01_n456 ) , .A2( us01_n507 ) , .A1( us01_n597 ) , .A4( us01_n626 ) , .A3( us01_n709 ) );
  NOR3_X1 us01_U9 (.A3( us01_n619 ) , .A2( us01_n620 ) , .ZN( us01_n634 ) , .A1( us01_n723 ) );
  NAND4_X1 us01_U90 (.A4( us01_n533 ) , .A3( us01_n534 ) , .A2( us01_n535 ) , .A1( us01_n536 ) , .ZN( us01_n620 ) );
  NOR4_X1 us01_U91 (.A4( us01_n524 ) , .A2( us01_n525 ) , .A1( us01_n526 ) , .ZN( us01_n536 ) , .A3( us01_n699 ) );
  NOR4_X1 us01_U92 (.A1( us01_n529 ) , .ZN( us01_n534 ) , .A2( us01_n652 ) , .A4( us01_n666 ) , .A3( us01_n763 ) );
  NOR4_X1 us01_U93 (.A4( us01_n527 ) , .A3( us01_n528 ) , .ZN( us01_n535 ) , .A2( us01_n682 ) , .A1( us01_n792 ) );
  NAND4_X1 us01_U94 (.A4( us01_n477 ) , .A3( us01_n478 ) , .A2( us01_n479 ) , .A1( us01_n480 ) , .ZN( us01_n692 ) );
  NOR3_X1 us01_U95 (.ZN( us01_n478 ) , .A2( us01_n506 ) , .A3( us01_n599 ) , .A1( us01_n608 ) );
  AOI211_X1 us01_U96 (.B( us01_n475 ) , .A( us01_n476 ) , .ZN( us01_n480 ) , .C2( us01_n831 ) , .C1( us01_n859 ) );
  NOR4_X1 us01_U97 (.ZN( us01_n479 ) , .A3( us01_n530 ) , .A4( us01_n543 ) , .A2( us01_n565 ) , .A1( us01_n715 ) );
  NAND4_X1 us01_U98 (.A4( us01_n546 ) , .A3( us01_n547 ) , .A2( us01_n548 ) , .A1( us01_n549 ) , .ZN( us01_n743 ) );
  NOR3_X1 us01_U99 (.ZN( us01_n547 ) , .A2( us01_n649 ) , .A1( us01_n665 ) , .A3( us01_n769 ) );
  NOR2_X1 us02_U10 (.ZN( us02_n574 ) , .A1( us02_n621 ) , .A2( us02_n744 ) );
  NOR2_X1 us02_U100 (.ZN( us02_n685 ) , .A1( us02_n830 ) , .A2( us02_n831 ) );
  NOR4_X1 us02_U101 (.ZN( us02_n619 ) , .A1( us02_n655 ) , .A3( us02_n665 ) , .A4( us02_n681 ) , .A2( us02_n765 ) );
  NOR4_X1 us02_U102 (.A4( us02_n608 ) , .A3( us02_n609 ) , .A2( us02_n610 ) , .A1( us02_n611 ) , .ZN( us02_n618 ) );
  NOR4_X1 us02_U103 (.A4( us02_n613 ) , .A3( us02_n614 ) , .A2( us02_n615 ) , .A1( us02_n616 ) , .ZN( us02_n617 ) );
  NAND4_X1 us02_U104 (.A4( us02_n484 ) , .A3( us02_n485 ) , .A2( us02_n486 ) , .A1( us02_n487 ) , .ZN( us02_n777 ) );
  NOR4_X1 us02_U105 (.A4( us02_n483 ) , .ZN( us02_n486 ) , .A1( us02_n565 ) , .A2( us02_n580 ) , .A3( us02_n601 ) );
  NOR4_X1 us02_U106 (.ZN( us02_n485 ) , .A1( us02_n506 ) , .A2( us02_n518 ) , .A4( us02_n545 ) , .A3( us02_n610 ) );
  NOR4_X1 us02_U107 (.ZN( us02_n484 ) , .A2( us02_n532 ) , .A1( us02_n557 ) , .A3( us02_n630 ) , .A4( us02_n717 ) );
  NAND4_X1 us02_U108 (.A4( us02_n690 ) , .A3( us02_n691 ) , .A1( us02_n692 ) , .ZN( us02_n775 ) , .A2( us02_n871 ) );
  AOI221_X1 us02_U109 (.A( us02_n680 ) , .ZN( us02_n691 ) , .B2( us02_n839 ) , .C1( us02_n841 ) , .C2( us02_n861 ) , .B1( us02_n864 ) );
  NOR2_X1 us02_U11 (.A1( us02_n677 ) , .ZN( us02_n692 ) , .A2( us02_n806 ) );
  INV_X1 us02_U110 (.A( us02_n678 ) , .ZN( us02_n871 ) );
  NOR4_X1 us02_U111 (.A4( us02_n686 ) , .A3( us02_n687 ) , .A2( us02_n688 ) , .A1( us02_n689 ) , .ZN( us02_n690 ) );
  NAND4_X1 us02_U112 (.A4( us02_n559 ) , .A3( us02_n560 ) , .A2( us02_n561 ) , .A1( us02_n562 ) , .ZN( us02_n606 ) );
  NOR4_X1 us02_U113 (.ZN( us02_n560 ) , .A1( us02_n652 ) , .A3( us02_n660 ) , .A4( us02_n684 ) , .A2( us02_n767 ) );
  NOR4_X1 us02_U114 (.A4( us02_n551 ) , .A3( us02_n552 ) , .A2( us02_n553 ) , .A1( us02_n554 ) , .ZN( us02_n561 ) );
  NOR4_X1 us02_U115 (.A4( us02_n555 ) , .A3( us02_n556 ) , .A2( us02_n557 ) , .A1( us02_n558 ) , .ZN( us02_n559 ) );
  NAND4_X1 us02_U116 (.A4( us02_n718 ) , .A3( us02_n719 ) , .A2( us02_n720 ) , .ZN( us02_n740 ) , .A1( us02_n856 ) );
  INV_X1 us02_U117 (.A( us02_n708 ) , .ZN( us02_n856 ) );
  AOI221_X1 us02_U118 (.A( us02_n709 ) , .ZN( us02_n720 ) , .C2( us02_n843 ) , .B2( us02_n844 ) , .C1( us02_n860 ) , .B1( us02_n861 ) );
  NOR4_X1 us02_U119 (.A4( us02_n714 ) , .A3( us02_n715 ) , .A2( us02_n716 ) , .A1( us02_n717 ) , .ZN( us02_n718 ) );
  INV_X1 us02_U12 (.A( us02_n679 ) , .ZN( us02_n839 ) );
  NAND4_X1 us02_U120 (.A4( us02_n472 ) , .A3( us02_n473 ) , .A2( us02_n474 ) , .A1( us02_n475 ) , .ZN( us02_n677 ) );
  NOR4_X1 us02_U121 (.A4( us02_n469 ) , .ZN( us02_n475 ) , .A3( us02_n555 ) , .A1( us02_n734 ) , .A2( us02_n754 ) );
  NOR4_X1 us02_U122 (.ZN( us02_n474 ) , .A1( us02_n530 ) , .A3( us02_n567 ) , .A4( us02_n599 ) , .A2( us02_n641 ) );
  NOR4_X1 us02_U123 (.ZN( us02_n473 ) , .A1( us02_n505 ) , .A3( us02_n543 ) , .A2( us02_n582 ) , .A4( us02_n715 ) );
  NOR2_X1 us02_U124 (.ZN( us02_n732 ) , .A2( us02_n831 ) , .A1( us02_n844 ) );
  NOR2_X1 us02_U125 (.ZN( us02_n788 ) , .A2( us02_n861 ) , .A1( us02_n867 ) );
  NOR2_X1 us02_U126 (.ZN( us02_n646 ) , .A1( us02_n853 ) , .A2( us02_n867 ) );
  NAND4_X1 us02_U127 (.A4( us02_n572 ) , .A3( us02_n573 ) , .A1( us02_n574 ) , .ZN( us02_n722 ) , .A2( us02_n873 ) );
  NOR4_X1 us02_U128 (.A4( us02_n568 ) , .A3( us02_n569 ) , .A2( us02_n570 ) , .A1( us02_n571 ) , .ZN( us02_n572 ) );
  AOI221_X1 us02_U129 (.A( us02_n563 ) , .C2( us02_n564 ) , .ZN( us02_n573 ) , .B2( us02_n844 ) , .B1( us02_n851 ) , .C1( us02_n852 ) );
  NOR4_X1 us02_U13 (.A4( us02_n444 ) , .A3( us02_n445 ) , .A2( us02_n515 ) , .A1( us02_n540 ) , .ZN( us02_n705 ) );
  INV_X1 us02_U130 (.A( us02_n606 ) , .ZN( us02_n873 ) );
  NAND4_X1 us02_U131 (.A4( us02_n492 ) , .A3( us02_n493 ) , .A1( us02_n494 ) , .ZN( us02_n801 ) , .A2( us02_n866 ) );
  AOI221_X1 us02_U132 (.A( us02_n488 ) , .ZN( us02_n493 ) , .B2( us02_n835 ) , .C2( us02_n840 ) , .C1( us02_n850 ) , .B1( us02_n859 ) );
  INV_X1 us02_U133 (.A( us02_n777 ) , .ZN( us02_n866 ) );
  NOR2_X1 us02_U134 (.ZN( us02_n494 ) , .A1( us02_n677 ) , .A2( us02_n693 ) );
  AOI222_X1 us02_U135 (.ZN( us02_n512 ) , .C1( us02_n831 ) , .B2( us02_n836 ) , .A2( us02_n842 ) , .C2( us02_n861 ) , .B1( us02_n862 ) , .A1( us02_n865 ) );
  NOR4_X1 us02_U136 (.A4( us02_n508 ) , .A2( us02_n509 ) , .A1( us02_n510 ) , .ZN( us02_n511 ) , .A3( us02_n669 ) );
  INV_X1 us02_U137 (.A( us02_n504 ) , .ZN( us02_n870 ) );
  INV_X1 us02_U138 (.A( us02_n761 ) , .ZN( us02_n829 ) );
  INV_X1 us02_U139 (.A( us02_n462 ) , .ZN( us02_n863 ) );
  OR3_X1 us02_U14 (.ZN( us02_n445 ) , .A1( us02_n527 ) , .A3( us02_n576 ) , .A2( us02_n874 ) );
  OAI21_X1 us02_U140 (.ZN( us02_n462 ) , .B1( us02_n808 ) , .A( us02_n833 ) , .B2( us02_n850 ) );
  OR4_X1 us02_U141 (.A4( us02_n565 ) , .A3( us02_n566 ) , .A2( us02_n567 ) , .ZN( us02_n571 ) , .A1( us02_n664 ) );
  OR4_X1 us02_U142 (.A4( us02_n517 ) , .A2( us02_n518 ) , .A1( us02_n519 ) , .ZN( us02_n521 ) , .A3( us02_n820 ) );
  OR4_X1 us02_U143 (.ZN( us02_n465 ) , .A4( us02_n517 ) , .A3( us02_n528 ) , .A2( us02_n577 ) , .A1( us02_n711 ) );
  OR4_X1 us02_U144 (.A4( us02_n681 ) , .A3( us02_n682 ) , .A2( us02_n683 ) , .A1( us02_n684 ) , .ZN( us02_n689 ) );
  OR4_X1 us02_U145 (.A4( us02_n579 ) , .A3( us02_n580 ) , .A2( us02_n581 ) , .A1( us02_n582 ) , .ZN( us02_n583 ) );
  NAND2_X1 us02_U146 (.ZN( us02_n612 ) , .A2( us02_n836 ) , .A1( us02_n872 ) );
  OR3_X1 us02_U147 (.A3( us02_n505 ) , .A2( us02_n506 ) , .A1( us02_n507 ) , .ZN( us02_n510 ) );
  AOI221_X1 us02_U148 (.A( us02_n712 ) , .B2( us02_n713 ) , .ZN( us02_n719 ) , .C1( us02_n831 ) , .B1( us02_n838 ) , .C2( us02_n862 ) );
  OR2_X1 us02_U149 (.A2( us02_n710 ) , .A1( us02_n711 ) , .ZN( us02_n712 ) );
  OR4_X1 us02_U15 (.A4( us02_n441 ) , .A2( us02_n442 ) , .A1( us02_n443 ) , .ZN( us02_n444 ) , .A3( us02_n552 ) );
  INV_X1 us02_U150 (.A( us02_n753 ) , .ZN( us02_n868 ) );
  OAI21_X1 us02_U151 (.B1( us02_n752 ) , .ZN( us02_n753 ) , .A( us02_n844 ) , .B2( us02_n867 ) );
  INV_X1 us02_U152 (.A( us02_n671 ) , .ZN( us02_n858 ) );
  AOI21_X1 us02_U153 (.A( us02_n669 ) , .B1( us02_n670 ) , .ZN( us02_n671 ) , .B2( us02_n855 ) );
  NAND2_X1 us02_U154 (.A1( us02_n446 ) , .A2( us02_n464 ) , .ZN( us02_n748 ) );
  OAI222_X1 us02_U155 (.B2( us02_n746 ) , .B1( us02_n747 ) , .A2( us02_n748 ) , .ZN( us02_n756 ) , .C2( us02_n804 ) , .C1( us02_n813 ) , .A1( us02_n816 ) );
  OAI222_X1 us02_U156 (.ZN( us02_n504 ) , .C2( us02_n624 ) , .B2( us02_n646 ) , .B1( us02_n746 ) , .A2( us02_n747 ) , .C1( us02_n804 ) , .A1( us02_n805 ) );
  OAI222_X1 us02_U157 (.B2( us02_n707 ) , .ZN( us02_n708 ) , .C2( us02_n723 ) , .B1( us02_n746 ) , .A1( us02_n805 ) , .C1( us02_n813 ) , .A2( us02_n814 ) );
  OAI222_X1 us02_U158 (.ZN( us02_n616 ) , .B1( us02_n696 ) , .C1( us02_n723 ) , .C2( us02_n746 ) , .B2( us02_n785 ) , .A2( us02_n791 ) , .A1( us02_n815 ) );
  NOR4_X1 us02_U159 (.A2( us02_n490 ) , .A1( us02_n491 ) , .ZN( us02_n492 ) , .A3( us02_n579 ) , .A4( us02_n611 ) );
  INV_X1 us02_U16 (.A( us02_n612 ) , .ZN( us02_n874 ) );
  OR4_X1 us02_U160 (.ZN( us02_n491 ) , .A4( us02_n533 ) , .A2( us02_n546 ) , .A1( us02_n558 ) , .A3( us02_n631 ) );
  OAI22_X1 us02_U161 (.B1( us02_n489 ) , .ZN( us02_n490 ) , .A1( us02_n685 ) , .A2( us02_n762 ) , .B2( us02_n816 ) );
  NOR3_X1 us02_U162 (.ZN( us02_n489 ) , .A1( us02_n781 ) , .A2( us02_n849 ) , .A3( us02_n862 ) );
  AOI22_X1 us02_U163 (.ZN( us02_n695 ) , .A1( us02_n829 ) , .B2( us02_n842 ) , .A2( us02_n864 ) , .B1( us02_n867 ) );
  INV_X1 us02_U164 (.A( us02_n729 ) , .ZN( us02_n838 ) );
  AOI221_X1 us02_U165 (.A( us02_n763 ) , .ZN( us02_n773 ) , .C2( us02_n809 ) , .B2( us02_n834 ) , .C1( us02_n854 ) , .B1( us02_n865 ) );
  AOI21_X1 us02_U166 (.B2( us02_n762 ) , .ZN( us02_n763 ) , .A( us02_n787 ) , .B1( us02_n791 ) );
  INV_X1 us02_U167 (.A( us02_n760 ) , .ZN( us02_n834 ) );
  AOI221_X1 us02_U168 (.A( us02_n482 ) , .ZN( us02_n487 ) , .B1( us02_n830 ) , .C2( us02_n843 ) , .C1( us02_n851 ) , .B2( us02_n861 ) );
  OAI22_X1 us02_U169 (.ZN( us02_n482 ) , .A1( us02_n707 ) , .B2( us02_n784 ) , .A2( us02_n805 ) , .B1( us02_n811 ) );
  INV_X1 us02_U17 (.A( us02_n748 ) , .ZN( us02_n862 ) );
  INV_X1 us02_U170 (.A( us02_n789 ) , .ZN( us02_n831 ) );
  NAND2_X1 us02_U171 (.A1( us02_n450 ) , .A2( us02_n452 ) , .ZN( us02_n761 ) );
  OAI221_X1 us02_U172 (.A( us02_n726 ) , .C2( us02_n727 ) , .B2( us02_n728 ) , .B1( us02_n729 ) , .ZN( us02_n736 ) , .C1( us02_n816 ) );
  AOI22_X1 us02_U173 (.ZN( us02_n726 ) , .B1( us02_n831 ) , .A2( us02_n837 ) , .A1( us02_n862 ) , .B2( us02_n865 ) );
  INV_X1 us02_U174 (.A( us02_n785 ) , .ZN( us02_n861 ) );
  OAI22_X1 us02_U175 (.ZN( us02_n709 ) , .A2( us02_n727 ) , .B2( us02_n728 ) , .A1( us02_n743 ) , .B1( us02_n812 ) );
  INV_X1 us02_U176 (.A( us02_n815 ) , .ZN( us02_n830 ) );
  OAI22_X1 us02_U177 (.ZN( us02_n488 ) , .A1( us02_n723 ) , .B2( us02_n727 ) , .B1( us02_n729 ) , .A2( us02_n778 ) );
  OAI22_X1 us02_U178 (.ZN( us02_n623 ) , .B1( us02_n668 ) , .B2( us02_n746 ) , .A1( us02_n814 ) , .A2( us02_n815 ) );
  INV_X1 us02_U179 (.A( us02_n743 ) , .ZN( us02_n836 ) );
  AOI222_X1 us02_U18 (.ZN( us02_n604 ) , .B2( us02_n670 ) , .B1( us02_n752 ) , .C2( us02_n830 ) , .A1( us02_n832 ) , .A2( us02_n861 ) , .C1( us02_n862 ) );
  OAI22_X1 us02_U180 (.A1( us02_n723 ) , .ZN( us02_n725 ) , .B2( us02_n749 ) , .B1( us02_n811 ) , .A2( us02_n815 ) );
  OAI22_X1 us02_U181 (.B2( us02_n778 ) , .B1( us02_n779 ) , .ZN( us02_n780 ) , .A2( us02_n813 ) , .A1( us02_n814 ) );
  INV_X1 us02_U182 (.A( us02_n787 ) , .ZN( us02_n844 ) );
  INV_X1 us02_U183 (.A( us02_n804 ) , .ZN( us02_n859 ) );
  INV_X1 us02_U184 (.A( us02_n813 ) , .ZN( us02_n832 ) );
  OAI22_X1 us02_U185 (.B2( us02_n743 ) , .ZN( us02_n745 ) , .A2( us02_n761 ) , .B1( us02_n779 ) , .A1( us02_n791 ) );
  OAI22_X1 us02_U186 (.B2( us02_n802 ) , .B1( us02_n803 ) , .A2( us02_n804 ) , .A1( us02_n805 ) , .ZN( us02_n807 ) );
  OAI22_X1 us02_U187 (.ZN( us02_n495 ) , .A2( us02_n743 ) , .A1( us02_n779 ) , .B1( us02_n790 ) , .B2( us02_n805 ) );
  OAI22_X1 us02_U188 (.ZN( us02_n589 ) , .B1( us02_n729 ) , .B2( us02_n748 ) , .A2( us02_n785 ) , .A1( us02_n802 ) );
  OAI22_X1 us02_U189 (.ZN( us02_n694 ) , .A2( us02_n729 ) , .A1( us02_n779 ) , .B1( us02_n790 ) , .B2( us02_n816 ) );
  AOI222_X1 us02_U19 (.ZN( us02_n562 ) , .B1( us02_n829 ) , .C1( us02_n840 ) , .A2( us02_n842 ) , .A1( us02_n853 ) , .B2( us02_n862 ) , .C2( us02_n872 ) );
  INV_X1 us02_U190 (.A( us02_n802 ) , .ZN( us02_n842 ) );
  INV_X1 us02_U191 (.A( us02_n668 ) , .ZN( us02_n864 ) );
  OAI22_X1 us02_U192 (.ZN( us02_n636 ) , .A1( us02_n698 ) , .B2( us02_n727 ) , .A2( us02_n761 ) , .B1( us02_n815 ) );
  NOR2_X1 us02_U193 (.ZN( us02_n714 ) , .A1( us02_n804 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U194 (.A1( us02_n696 ) , .ZN( us02_n769 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U195 (.ZN( us02_n665 ) , .A1( us02_n727 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U196 (.ZN( us02_n593 ) , .A2( us02_n696 ) , .A1( us02_n727 ) );
  NOR2_X1 us02_U197 (.ZN( us02_n569 ) , .A1( us02_n727 ) , .A2( us02_n805 ) );
  NOR2_X1 us02_U198 (.A2( us02_n743 ) , .ZN( us02_n754 ) , .A1( us02_n804 ) );
  NOR2_X1 us02_U199 (.ZN( us02_n717 ) , .A2( us02_n723 ) , .A1( us02_n743 ) );
  AOI222_X1 us02_U20 (.ZN( us02_n659 ) , .A2( us02_n838 ) , .B1( us02_n840 ) , .C2( us02_n844 ) , .A1( us02_n859 ) , .C1( us02_n862 ) , .B2( us02_n869 ) );
  NOR2_X1 us02_U200 (.ZN( us02_n734 ) , .A2( us02_n802 ) , .A1( us02_n804 ) );
  NOR2_X1 us02_U201 (.ZN( us02_n545 ) , .A2( us02_n779 ) , .A1( us02_n813 ) );
  NOR2_X1 us02_U202 (.ZN( us02_n576 ) , .A2( us02_n698 ) , .A1( us02_n813 ) );
  NOR2_X1 us02_U203 (.ZN( us02_n653 ) , .A1( us02_n727 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U204 (.ZN( us02_n611 ) , .A1( us02_n778 ) , .A2( us02_n785 ) );
  INV_X1 us02_U205 (.A( us02_n749 ) , .ZN( us02_n841 ) );
  NOR2_X1 us02_U206 (.ZN( us02_n531 ) , .A2( us02_n748 ) , .A1( us02_n749 ) );
  NOR2_X1 us02_U207 (.ZN( us02_n628 ) , .A2( us02_n727 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U208 (.ZN( us02_n614 ) , .A1( us02_n784 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U209 (.ZN( us02_n600 ) , .A2( us02_n779 ) , .A1( us02_n802 ) );
  INV_X1 us02_U21 (.A( us02_n646 ) , .ZN( us02_n869 ) );
  NOR2_X1 us02_U210 (.ZN( us02_n610 ) , .A2( us02_n779 ) , .A1( us02_n805 ) );
  INV_X1 us02_U211 (.A( us02_n746 ) , .ZN( us02_n833 ) );
  NOR2_X1 us02_U212 (.A2( us02_n743 ) , .ZN( us02_n768 ) , .A1( us02_n811 ) );
  NOR2_X1 us02_U213 (.ZN( us02_n527 ) , .A2( us02_n723 ) , .A1( us02_n802 ) );
  NOR2_X1 us02_U214 (.ZN( us02_n530 ) , .A2( us02_n779 ) , .A1( us02_n815 ) );
  NOR2_X1 us02_U215 (.ZN( us02_n627 ) , .A2( us02_n668 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U216 (.ZN( us02_n598 ) , .A2( us02_n790 ) , .A1( us02_n815 ) );
  INV_X1 us02_U217 (.A( us02_n727 ) , .ZN( us02_n851 ) );
  NOR2_X1 us02_U218 (.ZN( us02_n651 ) , .A1( us02_n668 ) , .A2( us02_n813 ) );
  NOR2_X1 us02_U219 (.A1( us02_n668 ) , .ZN( us02_n672 ) , .A2( us02_n743 ) );
  NOR4_X1 us02_U22 (.ZN( us02_n472 ) , .A2( us02_n520 ) , .A4( us02_n593 ) , .A1( us02_n608 ) , .A3( us02_n628 ) );
  NOR2_X1 us02_U220 (.ZN( us02_n601 ) , .A1( us02_n668 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U221 (.A1( us02_n668 ) , .ZN( us02_n687 ) , .A2( us02_n815 ) );
  INV_X1 us02_U222 (.A( us02_n791 ) , .ZN( us02_n850 ) );
  NOR2_X1 us02_U223 (.A2( us02_n707 ) , .A1( us02_n749 ) , .ZN( us02_n770 ) );
  NOR2_X1 us02_U224 (.A1( us02_n668 ) , .ZN( us02_n765 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U225 (.A1( us02_n698 ) , .ZN( us02_n767 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U226 (.ZN( us02_n540 ) , .A2( us02_n696 ) , .A1( us02_n698 ) );
  NOR2_X1 us02_U227 (.ZN( us02_n526 ) , .A1( us02_n668 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U228 (.ZN( us02_n666 ) , .A1( us02_n749 ) , .A2( us02_n814 ) );
  NOR2_X1 us02_U229 (.ZN( us02_n554 ) , .A1( us02_n749 ) , .A2( us02_n790 ) );
  NOR4_X1 us02_U23 (.ZN( us02_n478 ) , .A1( us02_n519 ) , .A4( us02_n556 ) , .A3( us02_n581 ) , .A2( us02_n629 ) );
  NOR2_X1 us02_U230 (.ZN( us02_n507 ) , .A2( us02_n779 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U231 (.ZN( us02_n542 ) , .A2( us02_n707 ) , .A1( us02_n784 ) );
  NOR2_X1 us02_U232 (.ZN( us02_n663 ) , .A1( us02_n784 ) , .A2( us02_n790 ) );
  NOR2_X1 us02_U233 (.A2( us02_n696 ) , .ZN( us02_n715 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U234 (.ZN( us02_n506 ) , .A1( us02_n811 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U235 (.ZN( us02_n555 ) , .A1( us02_n761 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U236 (.ZN( us02_n660 ) , .A1( us02_n728 ) , .A2( us02_n789 ) );
  NOR2_X1 us02_U237 (.ZN( us02_n661 ) , .A2( us02_n696 ) , .A1( us02_n728 ) );
  NOR2_X1 us02_U238 (.ZN( us02_n556 ) , .A1( us02_n791 ) , .A2( us02_n813 ) );
  NOR2_X1 us02_U239 (.ZN( us02_n544 ) , .A1( us02_n748 ) , .A2( us02_n813 ) );
  NOR4_X1 us02_U24 (.A4( us02_n531 ) , .A3( us02_n532 ) , .A2( us02_n533 ) , .ZN( us02_n534 ) , .A1( us02_n819 ) );
  NOR2_X1 us02_U240 (.ZN( us02_n508 ) , .A1( us02_n728 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U241 (.A2( us02_n696 ) , .A1( us02_n779 ) , .ZN( us02_n819 ) );
  OAI22_X1 us02_U242 (.B2( us02_n749 ) , .B1( us02_n750 ) , .A1( us02_n751 ) , .ZN( us02_n755 ) , .A2( us02_n805 ) );
  NOR2_X1 us02_U243 (.ZN( us02_n750 ) , .A2( us02_n851 ) , .A1( us02_n859 ) );
  NOR3_X1 us02_U244 (.ZN( us02_n751 ) , .A2( us02_n852 ) , .A1( us02_n862 ) , .A3( us02_n864 ) );
  NOR2_X1 us02_U245 (.ZN( us02_n529 ) , .A2( us02_n743 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U246 (.A1( us02_n748 ) , .ZN( us02_n766 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U247 (.ZN( us02_n543 ) , .A2( us02_n784 ) , .A1( us02_n791 ) );
  NOR2_X1 us02_U248 (.ZN( us02_n662 ) , .A1( us02_n728 ) , .A2( us02_n784 ) );
  NOR2_X1 us02_U249 (.ZN( us02_n630 ) , .A1( us02_n723 ) , .A2( us02_n812 ) );
  NOR4_X1 us02_U25 (.ZN( us02_n455 ) , .A2( us02_n516 ) , .A1( us02_n542 ) , .A3( us02_n578 ) , .A4( us02_n614 ) );
  NOR2_X1 us02_U250 (.ZN( us02_n613 ) , .A1( us02_n761 ) , .A2( us02_n811 ) );
  OAI22_X1 us02_U251 (.B1( us02_n439 ) , .ZN( us02_n443 ) , .A2( us02_n727 ) , .A1( us02_n743 ) , .B2( us02_n748 ) );
  NOR3_X1 us02_U252 (.ZN( us02_n439 ) , .A2( us02_n835 ) , .A3( us02_n836 ) , .A1( us02_n845 ) );
  NOR2_X1 us02_U253 (.ZN( us02_n505 ) , .A2( us02_n727 ) , .A1( us02_n761 ) );
  NOR2_X1 us02_U254 (.ZN( us02_n515 ) , .A1( us02_n707 ) , .A2( us02_n743 ) );
  NOR2_X1 us02_U255 (.ZN( us02_n716 ) , .A2( us02_n743 ) , .A1( us02_n785 ) );
  NOR2_X1 us02_U256 (.ZN( us02_n553 ) , .A1( us02_n785 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U257 (.ZN( us02_n516 ) , .A1( us02_n707 ) , .A2( us02_n802 ) );
  NOR2_X1 us02_U258 (.ZN( us02_n557 ) , .A1( us02_n707 ) , .A2( us02_n815 ) );
  NOR2_X1 us02_U259 (.ZN( us02_n669 ) , .A1( us02_n789 ) , .A2( us02_n804 ) );
  NOR4_X1 us02_U26 (.A4( us02_n540 ) , .A3( us02_n541 ) , .A2( us02_n542 ) , .ZN( us02_n549 ) , .A1( us02_n687 ) );
  NOR2_X1 us02_U260 (.ZN( us02_n520 ) , .A1( us02_n789 ) , .A2( us02_n811 ) );
  NOR2_X1 us02_U261 (.ZN( us02_n629 ) , .A1( us02_n746 ) , .A2( us02_n814 ) );
  INV_X1 us02_U262 (.A( us02_n805 ) , .ZN( us02_n840 ) );
  AOI21_X1 us02_U263 (.ZN( us02_n570 ) , .B2( us02_n696 ) , .B1( us02_n805 ) , .A( us02_n811 ) );
  NOR2_X1 us02_U264 (.ZN( us02_n654 ) , .A1( us02_n789 ) , .A2( us02_n814 ) );
  INV_X1 us02_U265 (.A( us02_n762 ) , .ZN( us02_n865 ) );
  AOI21_X1 us02_U266 (.ZN( us02_n551 ) , .B1( us02_n668 ) , .A( us02_n696 ) , .B2( us02_n804 ) );
  NOR2_X1 us02_U267 (.ZN( us02_n667 ) , .A2( us02_n707 ) , .A1( us02_n789 ) );
  NOR2_X1 us02_U268 (.ZN( us02_n655 ) , .A1( us02_n746 ) , .A2( us02_n779 ) );
  NOR2_X1 us02_U269 (.ZN( us02_n541 ) , .A1( us02_n761 ) , .A2( us02_n790 ) );
  NOR2_X1 us02_U27 (.ZN( us02_n679 ) , .A2( us02_n833 ) , .A1( us02_n838 ) );
  NOR2_X1 us02_U270 (.ZN( us02_n700 ) , .A2( us02_n785 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U271 (.ZN( us02_n608 ) , .A2( us02_n723 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U272 (.A1( us02_n729 ) , .ZN( us02_n764 ) , .A2( us02_n785 ) );
  AOI21_X1 us02_U273 (.A( us02_n814 ) , .B2( us02_n815 ) , .B1( us02_n816 ) , .ZN( us02_n817 ) );
  INV_X1 us02_U274 (.A( us02_n728 ) , .ZN( us02_n867 ) );
  NOR2_X1 us02_U275 (.ZN( us02_n578 ) , .A2( us02_n707 ) , .A1( us02_n729 ) );
  NOR2_X1 us02_U276 (.ZN( us02_n532 ) , .A2( us02_n723 ) , .A1( us02_n729 ) );
  AOI21_X1 us02_U277 (.B1( us02_n624 ) , .ZN( us02_n626 ) , .A( us02_n762 ) , .B2( us02_n813 ) );
  AOI21_X1 us02_U278 (.A( us02_n811 ) , .B2( us02_n812 ) , .B1( us02_n813 ) , .ZN( us02_n818 ) );
  AOI21_X1 us02_U279 (.ZN( us02_n514 ) , .A( us02_n728 ) , .B1( us02_n749 ) , .B2( us02_n802 ) );
  AOI222_X1 us02_U28 (.ZN( us02_n468 ) , .B1( us02_n831 ) , .A1( us02_n838 ) , .C1( us02_n841 ) , .C2( us02_n850 ) , .A2( us02_n854 ) , .B2( us02_n864 ) );
  AOI21_X1 us02_U280 (.ZN( us02_n498 ) , .B1( us02_n679 ) , .A( us02_n811 ) , .B2( us02_n815 ) );
  AOI21_X1 us02_U281 (.ZN( us02_n649 ) , .A( us02_n778 ) , .B1( us02_n791 ) , .B2( us02_n804 ) );
  AOI21_X1 us02_U282 (.ZN( us02_n477 ) , .B2( us02_n696 ) , .A( us02_n748 ) , .B1( us02_n778 ) );
  NOR2_X1 us02_U283 (.ZN( us02_n581 ) , .A1( us02_n743 ) , .A2( us02_n814 ) );
  AOI21_X1 us02_U284 (.ZN( us02_n592 ) , .B1( us02_n749 ) , .A( us02_n791 ) , .B2( us02_n812 ) );
  NOR2_X1 us02_U285 (.A2( us02_n707 ) , .A1( us02_n761 ) , .ZN( us02_n793 ) );
  AOI21_X1 us02_U286 (.ZN( us02_n625 ) , .B2( us02_n668 ) , .A( us02_n789 ) , .B1( us02_n790 ) );
  NOR2_X1 us02_U287 (.ZN( us02_n519 ) , .A2( us02_n707 ) , .A1( us02_n813 ) );
  AOI21_X1 us02_U288 (.ZN( us02_n476 ) , .A( us02_n668 ) , .B1( us02_n749 ) , .B2( us02_n805 ) );
  NOR2_X1 us02_U289 (.ZN( us02_n558 ) , .A2( us02_n790 ) , .A1( us02_n802 ) );
  NOR4_X1 us02_U29 (.A1( us02_n465 ) , .ZN( us02_n466 ) , .A4( us02_n541 ) , .A2( us02_n553 ) , .A3( us02_n613 ) );
  NOR2_X1 us02_U290 (.ZN( us02_n518 ) , .A2( us02_n698 ) , .A1( us02_n815 ) );
  NOR2_X1 us02_U291 (.ZN( us02_n682 ) , .A2( us02_n698 ) , .A1( us02_n802 ) );
  NOR2_X1 us02_U292 (.ZN( us02_n652 ) , .A1( us02_n761 ) , .A2( us02_n785 ) );
  INV_X1 us02_U293 (.A( us02_n812 ) , .ZN( us02_n835 ) );
  AOI21_X1 us02_U294 (.ZN( us02_n509 ) , .B2( us02_n668 ) , .A( us02_n729 ) , .B1( us02_n814 ) );
  AOI21_X1 us02_U295 (.ZN( us02_n538 ) , .B2( us02_n811 ) , .A( us02_n813 ) , .B1( us02_n814 ) );
  AOI21_X1 us02_U296 (.ZN( us02_n539 ) , .A( us02_n762 ) , .B2( us02_n778 ) , .B1( us02_n816 ) );
  NOR2_X1 us02_U297 (.ZN( us02_n580 ) , .A1( us02_n668 ) , .A2( us02_n787 ) );
  AOI21_X1 us02_U298 (.ZN( us02_n588 ) , .B2( us02_n698 ) , .B1( us02_n814 ) , .A( us02_n816 ) );
  AOI21_X1 us02_U299 (.B1( us02_n698 ) , .ZN( us02_n699 ) , .A( us02_n731 ) , .B2( us02_n762 ) );
  NAND2_X1 us02_U3 (.A1( us02_n440 ) , .A2( us02_n463 ) , .ZN( us02_n707 ) );
  AOI221_X1 us02_U30 (.ZN( us02_n467 ) , .C2( us02_n713 ) , .B2( us02_n830 ) , .C1( us02_n844 ) , .B1( us02_n859 ) , .A( us02_n863 ) );
  AOI21_X1 us02_U300 (.ZN( us02_n590 ) , .B2( us02_n762 ) , .A( us02_n784 ) , .B1( us02_n811 ) );
  AOI21_X1 us02_U301 (.ZN( us02_n497 ) , .A( us02_n723 ) , .B2( us02_n761 ) , .B1( us02_n813 ) );
  NOR2_X1 us02_U302 (.ZN( us02_n546 ) , .A1( us02_n698 ) , .A2( us02_n743 ) );
  INV_X1 us02_U303 (.A( us02_n790 ) , .ZN( us02_n872 ) );
  INV_X1 us02_U304 (.A( us02_n811 ) , .ZN( us02_n853 ) );
  AOI21_X1 us02_U305 (.ZN( us02_n648 ) , .B1( us02_n728 ) , .B2( us02_n762 ) , .A( us02_n812 ) );
  NOR2_X1 us02_U306 (.ZN( us02_n684 ) , .A1( us02_n728 ) , .A2( us02_n815 ) );
  AOI21_X1 us02_U307 (.B1( us02_n685 ) , .ZN( us02_n686 ) , .A( us02_n727 ) , .B2( us02_n760 ) );
  AOI21_X1 us02_U308 (.ZN( us02_n568 ) , .B1( us02_n749 ) , .B2( us02_n761 ) , .A( us02_n779 ) );
  AOI21_X1 us02_U309 (.ZN( us02_n499 ) , .A( us02_n696 ) , .B1( us02_n707 ) , .B2( us02_n785 ) );
  NOR4_X1 us02_U31 (.A4( us02_n513 ) , .A3( us02_n514 ) , .A2( us02_n515 ) , .A1( us02_n516 ) , .ZN( us02_n523 ) );
  NOR2_X1 us02_U310 (.ZN( us02_n567 ) , .A1( us02_n728 ) , .A2( us02_n761 ) );
  NOR2_X1 us02_U311 (.ZN( us02_n579 ) , .A2( us02_n696 ) , .A1( us02_n790 ) );
  NOR2_X1 us02_U312 (.ZN( us02_n565 ) , .A2( us02_n696 ) , .A1( us02_n762 ) );
  AOI21_X1 us02_U313 (.ZN( us02_n513 ) , .A( us02_n778 ) , .B2( us02_n791 ) , .B1( us02_n811 ) );
  INV_X1 us02_U314 (.A( us02_n698 ) , .ZN( us02_n852 ) );
  NOR2_X1 us02_U315 (.ZN( us02_n664 ) , .A1( us02_n779 ) , .A2( us02_n812 ) );
  AOI21_X1 us02_U316 (.ZN( us02_n449 ) , .B2( us02_n791 ) , .A( us02_n802 ) , .B1( us02_n814 ) );
  NOR2_X1 us02_U317 (.ZN( us02_n631 ) , .A2( us02_n696 ) , .A1( us02_n723 ) );
  AOI21_X1 us02_U318 (.ZN( us02_n563 ) , .B1( us02_n723 ) , .A( us02_n778 ) , .B2( us02_n790 ) );
  AOI21_X1 us02_U319 (.ZN( us02_n496 ) , .A( us02_n778 ) , .B2( us02_n790 ) , .B1( us02_n803 ) );
  AOI222_X1 us02_U32 (.ZN( us02_n524 ) , .A1( us02_n833 ) , .B2( us02_n836 ) , .C1( us02_n843 ) , .C2( us02_n849 ) , .A2( us02_n851 ) , .B1( us02_n865 ) );
  NAND2_X1 us02_U320 (.ZN( us02_n752 ) , .A1( us02_n762 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U321 (.ZN( us02_n528 ) , .A1( us02_n707 ) , .A2( us02_n778 ) );
  NOR2_X1 us02_U322 (.ZN( us02_n577 ) , .A1( us02_n707 ) , .A2( us02_n812 ) );
  AOI21_X1 us02_U323 (.ZN( us02_n688 ) , .B2( us02_n748 ) , .B1( us02_n762 ) , .A( us02_n805 ) );
  NOR2_X1 us02_U324 (.ZN( us02_n566 ) , .A1( us02_n746 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U325 (.ZN( us02_n683 ) , .A1( us02_n790 ) , .A2( us02_n812 ) );
  NOR2_X1 us02_U326 (.A2( us02_n812 ) , .A1( us02_n814 ) , .ZN( us02_n820 ) );
  AOI21_X1 us02_U327 (.A( us02_n789 ) , .B2( us02_n790 ) , .B1( us02_n791 ) , .ZN( us02_n792 ) );
  AOI21_X1 us02_U328 (.A( us02_n732 ) , .ZN( us02_n733 ) , .B2( us02_n779 ) , .B1( us02_n791 ) );
  NOR2_X1 us02_U329 (.ZN( us02_n710 ) , .A1( us02_n761 ) , .A2( us02_n762 ) );
  NOR4_X1 us02_U33 (.A3( us02_n520 ) , .A1( us02_n521 ) , .ZN( us02_n522 ) , .A2( us02_n672 ) , .A4( us02_n768 ) );
  NOR2_X1 us02_U330 (.ZN( us02_n582 ) , .A1( us02_n791 ) , .A2( us02_n816 ) );
  NOR2_X1 us02_U331 (.ZN( us02_n533 ) , .A1( us02_n723 ) , .A2( us02_n787 ) );
  NOR2_X1 us02_U332 (.ZN( us02_n681 ) , .A2( us02_n707 ) , .A1( us02_n816 ) );
  INV_X1 us02_U333 (.A( us02_n696 ) , .ZN( us02_n837 ) );
  NOR2_X1 us02_U334 (.ZN( us02_n641 ) , .A2( us02_n787 ) , .A1( us02_n790 ) );
  INV_X1 us02_U335 (.A( us02_n814 ) , .ZN( us02_n854 ) );
  AOI21_X1 us02_U336 (.ZN( us02_n441 ) , .A( us02_n698 ) , .B1( us02_n732 ) , .B2( us02_n749 ) );
  INV_X1 us02_U337 (.A( us02_n779 ) , .ZN( us02_n849 ) );
  AOI22_X1 us02_U338 (.A2( us02_n781 ) , .ZN( us02_n782 ) , .B2( us02_n830 ) , .A1( us02_n833 ) , .B1( us02_n862 ) );
  NAND2_X1 us02_U339 (.ZN( us02_n670 ) , .A1( us02_n805 ) , .A2( us02_n815 ) );
  NOR4_X1 us02_U34 (.A3( us02_n754 ) , .A2( us02_n755 ) , .A1( us02_n756 ) , .ZN( us02_n757 ) , .A4( us02_n868 ) );
  NAND2_X1 us02_U340 (.ZN( us02_n713 ) , .A1( us02_n727 ) , .A2( us02_n779 ) );
  NAND2_X1 us02_U341 (.A2( us02_n761 ) , .A1( us02_n805 ) , .ZN( us02_n809 ) );
  AOI21_X1 us02_U342 (.ZN( us02_n442 ) , .B1( us02_n788 ) , .B2( us02_n790 ) , .A( us02_n813 ) );
  NOR2_X1 us02_U343 (.ZN( us02_n483 ) , .A1( us02_n787 ) , .A2( us02_n804 ) );
  NOR2_X1 us02_U344 (.ZN( us02_n469 ) , .A2( us02_n778 ) , .A1( us02_n814 ) );
  INV_X1 us02_U345 (.A( us02_n784 ) , .ZN( us02_n845 ) );
  OAI21_X1 us02_U346 (.A( us02_n786 ) , .B2( us02_n787 ) , .B1( us02_n788 ) , .ZN( us02_n794 ) );
  OAI21_X1 us02_U347 (.ZN( us02_n786 ) , .A( us02_n838 ) , .B1( us02_n862 ) , .B2( us02_n872 ) );
  NOR2_X1 us02_U348 (.ZN( us02_n711 ) , .A2( us02_n723 ) , .A1( us02_n789 ) );
  NOR2_X1 us02_U349 (.ZN( us02_n525 ) , .A1( us02_n723 ) , .A2( us02_n749 ) );
  AOI211_X1 us02_U35 (.B( us02_n744 ) , .A( us02_n745 ) , .ZN( us02_n758 ) , .C1( us02_n831 ) , .C2( us02_n852 ) );
  NAND2_X1 us02_U350 (.A1( us02_n698 ) , .A2( us02_n728 ) , .ZN( us02_n781 ) );
  AOI21_X1 us02_U351 (.ZN( us02_n638 ) , .B2( us02_n748 ) , .A( us02_n787 ) , .B1( us02_n811 ) );
  AOI21_X1 us02_U352 (.ZN( us02_n639 ) , .B2( us02_n746 ) , .A( us02_n791 ) , .B1( us02_n802 ) );
  AOI21_X1 us02_U353 (.ZN( us02_n640 ) , .B1( us02_n679 ) , .A( us02_n790 ) , .B2( us02_n816 ) );
  NOR2_X1 us02_U354 (.ZN( us02_n517 ) , .A1( us02_n707 ) , .A2( us02_n787 ) );
  OAI21_X1 us02_U355 (.A( us02_n697 ) , .ZN( us02_n701 ) , .B2( us02_n749 ) , .B1( us02_n803 ) );
  OAI21_X1 us02_U356 (.ZN( us02_n697 ) , .B2( us02_n832 ) , .B1( us02_n837 ) , .A( us02_n859 ) );
  OAI21_X1 us02_U357 (.A( us02_n730 ) , .B1( us02_n731 ) , .ZN( us02_n735 ) , .B2( us02_n804 ) );
  OAI21_X1 us02_U358 (.ZN( us02_n730 ) , .A( us02_n832 ) , .B2( us02_n851 ) , .B1( us02_n872 ) );
  NAND2_X1 us02_U359 (.A2( us02_n748 ) , .A1( us02_n785 ) , .ZN( us02_n808 ) );
  NOR3_X1 us02_U36 (.A3( us02_n740 ) , .A2( us02_n741 ) , .A1( us02_n742 ) , .ZN( us02_n759 ) );
  INV_X1 us02_U360 (.A( us02_n816 ) , .ZN( us02_n843 ) );
  INV_X1 us02_U361 (.A( us02_n723 ) , .ZN( us02_n855 ) );
  AND2_X1 us02_U362 (.ZN( us02_n731 ) , .A1( us02_n778 ) , .A2( us02_n784 ) );
  NAND2_X1 us02_U363 (.A1( us02_n446 ) , .A2( us02_n448 ) , .ZN( us02_n804 ) );
  NAND2_X1 us02_U364 (.A1( us02_n454 ) , .A2( us02_n470 ) , .ZN( us02_n802 ) );
  NAND2_X1 us02_U365 (.A1( us02_n450 ) , .A2( us02_n453 ) , .ZN( us02_n813 ) );
  NAND2_X1 us02_U366 (.A1( us02_n450 ) , .A2( us02_n470 ) , .ZN( us02_n815 ) );
  NAND2_X1 us02_U367 (.A1( us02_n453 ) , .A2( us02_n460 ) , .ZN( us02_n812 ) );
  NAND2_X1 us02_U368 (.A1( us02_n452 ) , .A2( us02_n460 ) , .ZN( us02_n743 ) );
  NAND2_X1 us02_U369 (.A1( us02_n451 ) , .A2( us02_n464 ) , .ZN( us02_n668 ) );
  NOR4_X1 us02_U37 (.A4( us02_n733 ) , .A3( us02_n734 ) , .A2( us02_n735 ) , .A1( us02_n736 ) , .ZN( us02_n737 ) );
  NAND2_X1 us02_U370 (.A2( us02_n447 ) , .A1( us02_n459 ) , .ZN( us02_n727 ) );
  NAND2_X1 us02_U371 (.A1( us02_n454 ) , .A2( us02_n461 ) , .ZN( us02_n749 ) );
  NAND2_X1 us02_U372 (.A2( us02_n452 ) , .A1( us02_n454 ) , .ZN( us02_n805 ) );
  NAND2_X1 us02_U373 (.A2( us02_n453 ) , .A1( us02_n471 ) , .ZN( us02_n778 ) );
  NAND2_X1 us02_U374 (.A1( us02_n452 ) , .A2( us02_n471 ) , .ZN( us02_n784 ) );
  NAND2_X1 us02_U375 (.A2( us02_n463 ) , .A1( us02_n464 ) , .ZN( us02_n811 ) );
  NAND2_X1 us02_U376 (.A1( us02_n440 ) , .A2( us02_n459 ) , .ZN( us02_n698 ) );
  NAND2_X1 us02_U377 (.A2( us02_n448 ) , .A1( us02_n451 ) , .ZN( us02_n762 ) );
  NAND2_X1 us02_U378 (.A2( us02_n447 ) , .A1( us02_n451 ) , .ZN( us02_n728 ) );
  NAND2_X1 us02_U379 (.A2( us02_n460 ) , .A1( us02_n461 ) , .ZN( us02_n746 ) );
  AOI211_X1 us02_U38 (.B( us02_n724 ) , .A( us02_n725 ) , .ZN( us02_n738 ) , .C1( us02_n842 ) , .C2( us02_n854 ) );
  NAND2_X2 us02_U380 (.A2( us02_n460 ) , .A1( us02_n470 ) , .ZN( us02_n696 ) );
  NAND2_X1 us02_U381 (.A1( us02_n461 ) , .A2( us02_n471 ) , .ZN( us02_n787 ) );
  NOR2_X1 us02_U382 (.ZN( us02_n464 ) , .A2( us02_n846 ) , .A1( us02_n847 ) );
  NOR2_X1 us02_U383 (.ZN( us02_n452 ) , .A1( us02_n825 ) , .A2( us02_n826 ) );
  NOR2_X1 us02_U384 (.ZN( us02_n450 ) , .A1( us02_n827 ) , .A2( us02_n828 ) );
  NOR2_X1 us02_U385 (.ZN( us02_n446 ) , .A2( us02_n848 ) , .A1( us02_n857 ) );
  NAND2_X1 us02_U386 (.A2( us02_n453 ) , .A1( us02_n454 ) , .ZN( us02_n729 ) );
  NAND2_X1 us02_U387 (.A1( us02_n450 ) , .A2( us02_n461 ) , .ZN( us02_n789 ) );
  NAND2_X2 us02_U388 (.A2( us02_n447 ) , .A1( us02_n463 ) , .ZN( us02_n814 ) );
  NAND2_X2 us02_U389 (.A2( us02_n440 ) , .A1( us02_n451 ) , .ZN( us02_n790 ) );
  NOR3_X1 us02_U39 (.A3( us02_n721 ) , .A1( us02_n722 ) , .ZN( us02_n739 ) , .A2( us02_n740 ) );
  NAND2_X2 us02_U390 (.A1( us02_n448 ) , .A2( us02_n463 ) , .ZN( us02_n723 ) );
  NAND2_X1 us02_U391 (.A2( us02_n440 ) , .A1( us02_n446 ) , .ZN( us02_n783 ) );
  NAND2_X2 us02_U392 (.A1( us02_n448 ) , .A2( us02_n459 ) , .ZN( us02_n791 ) );
  NAND2_X2 us02_U393 (.A2( us02_n459 ) , .A1( us02_n464 ) , .ZN( us02_n779 ) );
  NAND2_X1 us02_U394 (.A1( us02_n446 ) , .A2( us02_n447 ) , .ZN( us02_n785 ) );
  NOR2_X1 us02_U395 (.A2( sa02_6 ) , .A1( sa02_7 ) , .ZN( us02_n463 ) );
  NOR2_X1 us02_U396 (.A2( sa02_5 ) , .ZN( us02_n447 ) , .A1( us02_n846 ) );
  NOR2_X1 us02_U397 (.A2( sa02_7 ) , .ZN( us02_n459 ) , .A1( us02_n848 ) );
  NOR2_X1 us02_U398 (.A2( sa02_4 ) , .ZN( us02_n448 ) , .A1( us02_n847 ) );
  NOR2_X1 us02_U399 (.A2( sa02_4 ) , .A1( sa02_5 ) , .ZN( us02_n440 ) );
  NAND2_X1 us02_U4 (.A2( us02_n470 ) , .A1( us02_n471 ) , .ZN( us02_n816 ) );
  AOI221_X1 us02_U40 (.A( us02_n780 ) , .ZN( us02_n797 ) , .C2( us02_n836 ) , .B2( us02_n837 ) , .B1( us02_n864 ) , .C1( us02_n865 ) );
  NOR2_X1 us02_U400 (.A2( sa02_1 ) , .ZN( us02_n470 ) , .A1( us02_n825 ) );
  NOR2_X1 us02_U401 (.A2( sa02_2 ) , .A1( sa02_3 ) , .ZN( us02_n471 ) );
  NOR2_X1 us02_U402 (.A2( sa02_6 ) , .ZN( us02_n451 ) , .A1( us02_n857 ) );
  NOR2_X1 us02_U403 (.A2( sa02_2 ) , .ZN( us02_n460 ) , .A1( us02_n828 ) );
  NOR2_X1 us02_U404 (.A2( sa02_0 ) , .ZN( us02_n453 ) , .A1( us02_n826 ) );
  NOR2_X1 us02_U405 (.A2( sa02_0 ) , .A1( sa02_1 ) , .ZN( us02_n461 ) );
  NOR2_X1 us02_U406 (.A2( sa02_3 ) , .ZN( us02_n454 ) , .A1( us02_n827 ) );
  INV_X1 us02_U407 (.A( sa02_6 ) , .ZN( us02_n848 ) );
  INV_X1 us02_U408 (.A( sa02_1 ) , .ZN( us02_n826 ) );
  INV_X1 us02_U409 (.A( sa02_3 ) , .ZN( us02_n828 ) );
  NOR4_X1 us02_U41 (.A4( us02_n792 ) , .A3( us02_n793 ) , .A2( us02_n794 ) , .A1( us02_n795 ) , .ZN( us02_n796 ) );
  INV_X1 us02_U410 (.A( sa02_2 ) , .ZN( us02_n827 ) );
  INV_X1 us02_U411 (.A( sa02_0 ) , .ZN( us02_n825 ) );
  INV_X1 us02_U412 (.A( sa02_5 ) , .ZN( us02_n847 ) );
  INV_X1 us02_U413 (.A( sa02_7 ) , .ZN( us02_n857 ) );
  OAI221_X1 us02_U414 (.A( us02_n782 ) , .C2( us02_n783 ) , .B2( us02_n784 ) , .B1( us02_n785 ) , .ZN( us02_n795 ) , .C1( us02_n812 ) );
  OAI22_X1 us02_U415 (.ZN( us02_n587 ) , .A2( us02_n746 ) , .B2( us02_n761 ) , .A1( us02_n762 ) , .B1( us02_n783 ) );
  AOI21_X1 us02_U416 (.ZN( us02_n591 ) , .B1( us02_n727 ) , .B2( us02_n783 ) , .A( us02_n789 ) );
  OAI221_X1 us02_U417 (.A( us02_n695 ) , .ZN( us02_n702 ) , .C2( us02_n783 ) , .C1( us02_n784 ) , .B1( us02_n785 ) , .B2( us02_n805 ) );
  NAND2_X1 us02_U418 (.A1( us02_n728 ) , .A2( us02_n783 ) , .ZN( us02_n810 ) );
  AOI21_X1 us02_U419 (.ZN( us02_n622 ) , .B1( us02_n698 ) , .A( us02_n778 ) , .B2( us02_n783 ) );
  NOR4_X1 us02_U42 (.A4( us02_n775 ) , .A3( us02_n776 ) , .A1( us02_n777 ) , .ZN( us02_n798 ) , .A2( us02_n800 ) );
  OAI22_X1 us02_U420 (.ZN( us02_n680 ) , .A1( us02_n698 ) , .A2( us02_n729 ) , .B2( us02_n783 ) , .B1( us02_n816 ) );
  AOI21_X1 us02_U421 (.ZN( us02_n647 ) , .A( us02_n761 ) , .B2( us02_n783 ) , .B1( us02_n791 ) );
  OAI21_X1 us02_U422 (.A( us02_n612 ) , .ZN( us02_n615 ) , .B1( us02_n624 ) , .B2( us02_n783 ) );
  NOR2_X1 us02_U423 (.ZN( us02_n650 ) , .A1( us02_n783 ) , .A2( us02_n787 ) );
  NOR2_X1 us02_U424 (.ZN( us02_n552 ) , .A2( us02_n743 ) , .A1( us02_n783 ) );
  NOR2_X1 us02_U425 (.ZN( us02_n609 ) , .A1( us02_n783 ) , .A2( us02_n815 ) );
  OAI222_X1 us02_U426 (.A2( us02_n668 ) , .ZN( us02_n673 ) , .B1( us02_n746 ) , .B2( us02_n783 ) , .C2( us02_n787 ) , .C1( us02_n814 ) , .A1( us02_n816 ) );
  NOR2_X1 us02_U427 (.ZN( us02_n599 ) , .A2( us02_n696 ) , .A1( us02_n783 ) );
  INV_X1 us02_U428 (.A( us02_n783 ) , .ZN( us02_n860 ) );
  AOI221_X1 us02_U429 (.A( us02_n575 ) , .ZN( us02_n586 ) , .B2( us02_n830 ) , .C2( us02_n842 ) , .B1( us02_n853 ) , .C1( us02_n860 ) );
  NOR2_X1 us02_U43 (.ZN( us02_n803 ) , .A1( us02_n853 ) , .A2( us02_n860 ) );
  AOI21_X1 us02_U430 (.ZN( us02_n575 ) , .B2( us02_n723 ) , .B1( us02_n747 ) , .A( us02_n784 ) );
  INV_X1 us02_U431 (.A( sa02_4 ) , .ZN( us02_n846 ) );
  NAND2_X1 us02_U432 (.ZN( sa02_sr_2 ) , .A2( us02_n438 ) , .A1( us02_n644 ) );
  NOR3_X1 us02_U433 (.A2( us02_n606 ) , .A1( us02_n607 ) , .ZN( us02_n645 ) , .A3( us02_n721 ) );
  AOI222_X1 us02_U434 (.B2( us02_n637 ) , .ZN( us02_n643 ) , .B1( us02_n840 ) , .A1( us02_n841 ) , .C2( us02_n845 ) , .C1( us02_n862 ) , .A2( us02_n864 ) );
  NOR4_X1 us02_U435 (.A4( us02_n638 ) , .A3( us02_n639 ) , .A2( us02_n640 ) , .A1( us02_n641 ) , .ZN( us02_n642 ) );
  AOI211_X1 us02_U436 (.A( us02_n636 ) , .ZN( us02_n644 ) , .B( us02_n742 ) , .C2( us02_n838 ) , .C1( us02_n853 ) );
  NAND3_X1 us02_U437 (.ZN( sa02_sr_6 ) , .A3( us02_n796 ) , .A2( us02_n797 ) , .A1( us02_n798 ) );
  NAND3_X1 us02_U438 (.ZN( sa02_sr_5 ) , .A3( us02_n757 ) , .A2( us02_n758 ) , .A1( us02_n759 ) );
  NAND3_X1 us02_U439 (.ZN( sa02_sr_4 ) , .A3( us02_n737 ) , .A2( us02_n738 ) , .A1( us02_n739 ) );
  NAND4_X1 us02_U44 (.ZN( sa02_sr_3 ) , .A4( us02_n703 ) , .A3( us02_n704 ) , .A2( us02_n705 ) , .A1( us02_n706 ) );
  NAND3_X1 us02_U440 (.A3( us02_n674 ) , .A2( us02_n675 ) , .A1( us02_n676 ) , .ZN( us02_n806 ) );
  NAND3_X1 us02_U441 (.ZN( us02_n637 ) , .A3( us02_n707 ) , .A2( us02_n723 ) , .A1( us02_n791 ) );
  NAND3_X1 us02_U442 (.A3( us02_n617 ) , .A2( us02_n618 ) , .A1( us02_n619 ) , .ZN( us02_n724 ) );
  NAND3_X1 us02_U443 (.A3( us02_n584 ) , .A2( us02_n585 ) , .A1( us02_n586 ) , .ZN( us02_n620 ) );
  NAND3_X1 us02_U444 (.ZN( us02_n564 ) , .A3( us02_n679 ) , .A2( us02_n749 ) , .A1( us02_n784 ) );
  NAND3_X1 us02_U445 (.A3( us02_n522 ) , .A2( us02_n523 ) , .A1( us02_n524 ) , .ZN( us02_n741 ) );
  NAND3_X1 us02_U446 (.A3( us02_n511 ) , .A1( us02_n512 ) , .ZN( us02_n607 ) , .A2( us02_n870 ) );
  NAND3_X1 us02_U447 (.A3( us02_n466 ) , .A2( us02_n467 ) , .A1( us02_n468 ) , .ZN( us02_n776 ) );
  NAND4_X1 us02_U448 (.A4( us02_n632 ) , .A3( us02_n633 ) , .A2( us02_n634 ) , .A1( us02_n635 ) , .ZN( us02_n742 ) );
  NOR4_X1 us02_U45 (.A4( us02_n699 ) , .A3( us02_n700 ) , .A2( us02_n701 ) , .A1( us02_n702 ) , .ZN( us02_n703 ) );
  AOI211_X1 us02_U46 (.B( us02_n693 ) , .A( us02_n694 ) , .ZN( us02_n704 ) , .C2( us02_n830 ) , .C1( us02_n850 ) );
  NOR2_X1 us02_U47 (.ZN( us02_n706 ) , .A2( us02_n775 ) , .A1( us02_n799 ) );
  NAND4_X1 us02_U48 (.ZN( sa02_sr_7 ) , .A4( us02_n821 ) , .A3( us02_n822 ) , .A2( us02_n823 ) , .A1( us02_n824 ) );
  NOR4_X1 us02_U49 (.A4( us02_n817 ) , .A3( us02_n818 ) , .A2( us02_n819 ) , .A1( us02_n820 ) , .ZN( us02_n821 ) );
  NOR3_X1 us02_U5 (.ZN( us02_n597 ) , .A1( us02_n607 ) , .A3( us02_n722 ) , .A2( us02_n741 ) );
  AOI222_X1 us02_U50 (.C2( us02_n808 ) , .B2( us02_n809 ) , .A2( us02_n810 ) , .ZN( us02_n822 ) , .C1( us02_n831 ) , .A1( us02_n838 ) , .B1( us02_n852 ) );
  AOI211_X1 us02_U51 (.B( us02_n806 ) , .A( us02_n807 ) , .ZN( us02_n823 ) , .C1( us02_n841 ) , .C2( us02_n849 ) );
  NOR2_X1 us02_U52 (.ZN( us02_n747 ) , .A1( us02_n860 ) , .A2( us02_n861 ) );
  NAND4_X1 us02_U53 (.ZN( sa02_sr_0 ) , .A4( us02_n500 ) , .A3( us02_n501 ) , .A2( us02_n502 ) , .A1( us02_n503 ) );
  AOI221_X1 us02_U54 (.A( us02_n496 ) , .ZN( us02_n501 ) , .B2( us02_n842 ) , .C1( us02_n845 ) , .C2( us02_n859 ) , .B1( us02_n861 ) );
  NOR4_X1 us02_U55 (.A4( us02_n497 ) , .A3( us02_n498 ) , .A2( us02_n499 ) , .ZN( us02_n500 ) , .A1( us02_n526 ) );
  AOI211_X1 us02_U56 (.A( us02_n495 ) , .ZN( us02_n502 ) , .B( us02_n801 ) , .C2( us02_n838 ) , .C1( us02_n850 ) );
  NAND4_X1 us02_U57 (.ZN( sa02_sr_1 ) , .A4( us02_n594 ) , .A3( us02_n595 ) , .A2( us02_n596 ) , .A1( us02_n597 ) );
  NOR4_X1 us02_U58 (.A4( us02_n590 ) , .A3( us02_n591 ) , .A2( us02_n592 ) , .A1( us02_n593 ) , .ZN( us02_n594 ) );
  AOI211_X1 us02_U59 (.B( us02_n588 ) , .A( us02_n589 ) , .ZN( us02_n595 ) , .C2( us02_n810 ) , .C1( us02_n832 ) );
  NOR3_X1 us02_U6 (.A3( us02_n799 ) , .A2( us02_n800 ) , .A1( us02_n801 ) , .ZN( us02_n824 ) );
  AOI211_X1 us02_U60 (.A( us02_n587 ) , .ZN( us02_n596 ) , .B( us02_n620 ) , .C1( us02_n844 ) , .C2( us02_n854 ) );
  NOR2_X1 us02_U61 (.ZN( us02_n624 ) , .A2( us02_n835 ) , .A1( us02_n838 ) );
  AND3_X1 us02_U62 (.ZN( us02_n438 ) , .A2( us02_n642 ) , .A3( us02_n643 ) , .A1( us02_n645 ) );
  NOR4_X1 us02_U63 (.A4( us02_n576 ) , .A3( us02_n577 ) , .A2( us02_n578 ) , .ZN( us02_n585 ) , .A1( us02_n682 ) );
  NOR4_X1 us02_U64 (.A1( us02_n583 ) , .ZN( us02_n584 ) , .A3( us02_n651 ) , .A2( us02_n661 ) , .A4( us02_n766 ) );
  AOI211_X1 us02_U65 (.B( us02_n622 ) , .A( us02_n623 ) , .ZN( us02_n634 ) , .C2( us02_n835 ) , .C1( us02_n862 ) );
  NOR4_X1 us02_U66 (.A4( us02_n628 ) , .A3( us02_n629 ) , .A2( us02_n630 ) , .A1( us02_n631 ) , .ZN( us02_n632 ) );
  NOR4_X1 us02_U67 (.A4( us02_n625 ) , .A3( us02_n626 ) , .A2( us02_n627 ) , .ZN( us02_n633 ) , .A1( us02_n663 ) );
  NAND4_X1 us02_U68 (.A4( us02_n656 ) , .A3( us02_n657 ) , .A2( us02_n658 ) , .A1( us02_n659 ) , .ZN( us02_n799 ) );
  NOR3_X1 us02_U69 (.A3( us02_n647 ) , .A2( us02_n648 ) , .A1( us02_n649 ) , .ZN( us02_n658 ) );
  NOR3_X1 us02_U7 (.ZN( us02_n503 ) , .A2( us02_n678 ) , .A3( us02_n776 ) , .A1( us02_n875 ) );
  NOR3_X1 us02_U70 (.A3( us02_n650 ) , .A2( us02_n651 ) , .A1( us02_n652 ) , .ZN( us02_n657 ) );
  NOR3_X1 us02_U71 (.A3( us02_n653 ) , .A2( us02_n654 ) , .A1( us02_n655 ) , .ZN( us02_n656 ) );
  NAND4_X1 us02_U72 (.A4( us02_n771 ) , .A3( us02_n772 ) , .A2( us02_n773 ) , .A1( us02_n774 ) , .ZN( us02_n800 ) );
  NOR3_X1 us02_U73 (.A3( us02_n764 ) , .A2( us02_n765 ) , .A1( us02_n766 ) , .ZN( us02_n772 ) );
  NOR4_X1 us02_U74 (.A4( us02_n767 ) , .A3( us02_n768 ) , .A2( us02_n769 ) , .A1( us02_n770 ) , .ZN( us02_n771 ) );
  AOI222_X1 us02_U75 (.ZN( us02_n774 ) , .A1( us02_n829 ) , .C1( us02_n833 ) , .B2( us02_n840 ) , .A2( us02_n849 ) , .B1( us02_n860 ) , .C2( us02_n872 ) );
  NOR4_X1 us02_U76 (.A4( us02_n664 ) , .A3( us02_n665 ) , .A2( us02_n666 ) , .A1( us02_n667 ) , .ZN( us02_n675 ) );
  NOR4_X1 us02_U77 (.A4( us02_n660 ) , .A3( us02_n661 ) , .A2( us02_n662 ) , .A1( us02_n663 ) , .ZN( us02_n676 ) );
  NOR4_X1 us02_U78 (.A3( us02_n672 ) , .A1( us02_n673 ) , .ZN( us02_n674 ) , .A4( us02_n714 ) , .A2( us02_n858 ) );
  NOR2_X1 us02_U79 (.ZN( us02_n760 ) , .A1( us02_n832 ) , .A2( us02_n833 ) );
  INV_X1 us02_U8 (.A( us02_n705 ) , .ZN( us02_n875 ) );
  NAND4_X1 us02_U80 (.A4( us02_n455 ) , .A3( us02_n456 ) , .A2( us02_n457 ) , .A1( us02_n458 ) , .ZN( us02_n678 ) );
  NOR3_X1 us02_U81 (.ZN( us02_n456 ) , .A3( us02_n529 ) , .A1( us02_n554 ) , .A2( us02_n569 ) );
  AOI221_X1 us02_U82 (.A( us02_n449 ) , .ZN( us02_n458 ) , .C2( us02_n752 ) , .B1( us02_n831 ) , .C1( us02_n841 ) , .B2( us02_n860 ) );
  NOR4_X1 us02_U83 (.ZN( us02_n457 ) , .A2( us02_n508 ) , .A1( us02_n598 ) , .A4( us02_n627 ) , .A3( us02_n710 ) );
  NAND4_X1 us02_U84 (.A4( us02_n602 ) , .A3( us02_n603 ) , .A2( us02_n604 ) , .A1( us02_n605 ) , .ZN( us02_n721 ) );
  NOR3_X1 us02_U85 (.A1( us02_n598 ) , .ZN( us02_n603 ) , .A3( us02_n662 ) , .A2( us02_n769 ) );
  NOR4_X1 us02_U86 (.A3( us02_n599 ) , .A2( us02_n600 ) , .A1( us02_n601 ) , .ZN( us02_n602 ) , .A4( us02_n654 ) );
  AOI222_X1 us02_U87 (.ZN( us02_n605 ) , .A1( us02_n829 ) , .C2( us02_n836 ) , .B1( us02_n841 ) , .A2( us02_n855 ) , .B2( us02_n860 ) , .C1( us02_n867 ) );
  NAND4_X1 us02_U88 (.A4( us02_n534 ) , .A3( us02_n535 ) , .A2( us02_n536 ) , .A1( us02_n537 ) , .ZN( us02_n621 ) );
  NOR4_X1 us02_U89 (.A4( us02_n525 ) , .A2( us02_n526 ) , .A1( us02_n527 ) , .ZN( us02_n537 ) , .A3( us02_n700 ) );
  NOR3_X1 us02_U9 (.A3( us02_n620 ) , .A2( us02_n621 ) , .ZN( us02_n635 ) , .A1( us02_n724 ) );
  NOR4_X1 us02_U90 (.A1( us02_n530 ) , .ZN( us02_n535 ) , .A2( us02_n653 ) , .A4( us02_n667 ) , .A3( us02_n764 ) );
  NOR4_X1 us02_U91 (.A4( us02_n528 ) , .A3( us02_n529 ) , .ZN( us02_n536 ) , .A2( us02_n683 ) , .A1( us02_n793 ) );
  NAND4_X1 us02_U92 (.A4( us02_n547 ) , .A3( us02_n548 ) , .A2( us02_n549 ) , .A1( us02_n550 ) , .ZN( us02_n744 ) );
  NOR3_X1 us02_U93 (.ZN( us02_n548 ) , .A2( us02_n650 ) , .A1( us02_n666 ) , .A3( us02_n770 ) );
  AOI211_X1 us02_U94 (.B( us02_n538 ) , .A( us02_n539 ) , .ZN( us02_n550 ) , .C2( us02_n838 ) , .C1( us02_n850 ) );
  NOR4_X1 us02_U95 (.A4( us02_n543 ) , .A3( us02_n544 ) , .A2( us02_n545 ) , .A1( us02_n546 ) , .ZN( us02_n547 ) );
  NAND4_X1 us02_U96 (.A4( us02_n478 ) , .A3( us02_n479 ) , .A2( us02_n480 ) , .A1( us02_n481 ) , .ZN( us02_n693 ) );
  NOR3_X1 us02_U97 (.ZN( us02_n479 ) , .A2( us02_n507 ) , .A3( us02_n600 ) , .A1( us02_n609 ) );
  AOI211_X1 us02_U98 (.B( us02_n476 ) , .A( us02_n477 ) , .ZN( us02_n481 ) , .C2( us02_n832 ) , .C1( us02_n860 ) );
  NOR4_X1 us02_U99 (.ZN( us02_n480 ) , .A3( us02_n531 ) , .A4( us02_n544 ) , .A2( us02_n566 ) , .A1( us02_n716 ) );
  NOR3_X1 us12_U10 (.ZN( us12_n504 ) , .A2( us12_n679 ) , .A3( us12_n777 ) , .A1( us12_n876 ) );
  NOR4_X1 us12_U100 (.A4( us12_n529 ) , .A3( us12_n530 ) , .ZN( us12_n537 ) , .A2( us12_n684 ) , .A1( us12_n794 ) );
  NAND4_X1 us12_U101 (.A4( us12_n479 ) , .A3( us12_n480 ) , .A2( us12_n481 ) , .A1( us12_n482 ) , .ZN( us12_n694 ) );
  NOR3_X1 us12_U102 (.ZN( us12_n480 ) , .A2( us12_n508 ) , .A3( us12_n601 ) , .A1( us12_n610 ) );
  AOI211_X1 us12_U103 (.B( us12_n477 ) , .A( us12_n478 ) , .ZN( us12_n482 ) , .C2( us12_n833 ) , .C1( us12_n861 ) );
  NOR4_X1 us12_U104 (.ZN( us12_n481 ) , .A3( us12_n532 ) , .A4( us12_n545 ) , .A2( us12_n567 ) , .A1( us12_n717 ) );
  NAND4_X1 us12_U105 (.A4( us12_n548 ) , .A3( us12_n549 ) , .A2( us12_n550 ) , .A1( us12_n551 ) , .ZN( us12_n745 ) );
  NOR3_X1 us12_U106 (.ZN( us12_n549 ) , .A2( us12_n651 ) , .A1( us12_n667 ) , .A3( us12_n771 ) );
  AOI211_X1 us12_U107 (.B( us12_n539 ) , .A( us12_n540 ) , .ZN( us12_n551 ) , .C2( us12_n839 ) , .C1( us12_n851 ) );
  NOR4_X1 us12_U108 (.A4( us12_n541 ) , .A3( us12_n542 ) , .A2( us12_n543 ) , .ZN( us12_n550 ) , .A1( us12_n688 ) );
  NOR4_X1 us12_U109 (.ZN( us12_n620 ) , .A1( us12_n656 ) , .A3( us12_n666 ) , .A4( us12_n682 ) , .A2( us12_n766 ) );
  INV_X1 us12_U11 (.A( us12_n706 ) , .ZN( us12_n876 ) );
  NOR4_X1 us12_U110 (.A4( us12_n609 ) , .A3( us12_n610 ) , .A2( us12_n611 ) , .A1( us12_n612 ) , .ZN( us12_n619 ) );
  NOR4_X1 us12_U111 (.A4( us12_n614 ) , .A3( us12_n615 ) , .A2( us12_n616 ) , .A1( us12_n617 ) , .ZN( us12_n618 ) );
  NOR2_X1 us12_U112 (.ZN( us12_n686 ) , .A1( us12_n831 ) , .A2( us12_n832 ) );
  NAND4_X1 us12_U113 (.A4( us12_n485 ) , .A3( us12_n486 ) , .A2( us12_n487 ) , .A1( us12_n488 ) , .ZN( us12_n778 ) );
  NOR4_X1 us12_U114 (.A4( us12_n484 ) , .ZN( us12_n487 ) , .A1( us12_n566 ) , .A2( us12_n581 ) , .A3( us12_n602 ) );
  NOR4_X1 us12_U115 (.ZN( us12_n486 ) , .A1( us12_n507 ) , .A2( us12_n519 ) , .A4( us12_n546 ) , .A3( us12_n611 ) );
  NOR4_X1 us12_U116 (.ZN( us12_n485 ) , .A2( us12_n533 ) , .A1( us12_n558 ) , .A3( us12_n631 ) , .A4( us12_n718 ) );
  NAND4_X1 us12_U117 (.A4( us12_n691 ) , .A3( us12_n692 ) , .A1( us12_n693 ) , .ZN( us12_n776 ) , .A2( us12_n872 ) );
  AOI221_X1 us12_U118 (.A( us12_n681 ) , .ZN( us12_n692 ) , .B2( us12_n840 ) , .C1( us12_n842 ) , .C2( us12_n862 ) , .B1( us12_n865 ) );
  INV_X1 us12_U119 (.A( us12_n679 ) , .ZN( us12_n872 ) );
  NOR3_X1 us12_U12 (.A3( us12_n621 ) , .A2( us12_n622 ) , .ZN( us12_n636 ) , .A1( us12_n725 ) );
  NOR4_X1 us12_U120 (.A4( us12_n687 ) , .A3( us12_n688 ) , .A2( us12_n689 ) , .A1( us12_n690 ) , .ZN( us12_n691 ) );
  NAND4_X1 us12_U121 (.A4( us12_n719 ) , .A3( us12_n720 ) , .A2( us12_n721 ) , .ZN( us12_n741 ) , .A1( us12_n857 ) );
  INV_X1 us12_U122 (.A( us12_n709 ) , .ZN( us12_n857 ) );
  AOI221_X1 us12_U123 (.A( us12_n710 ) , .ZN( us12_n721 ) , .C2( us12_n844 ) , .B2( us12_n845 ) , .C1( us12_n861 ) , .B1( us12_n862 ) );
  NOR4_X1 us12_U124 (.A4( us12_n715 ) , .A3( us12_n716 ) , .A2( us12_n717 ) , .A1( us12_n718 ) , .ZN( us12_n719 ) );
  NAND4_X1 us12_U125 (.A4( us12_n473 ) , .A3( us12_n474 ) , .A2( us12_n475 ) , .A1( us12_n476 ) , .ZN( us12_n678 ) );
  NOR4_X1 us12_U126 (.ZN( us12_n475 ) , .A1( us12_n531 ) , .A3( us12_n568 ) , .A4( us12_n600 ) , .A2( us12_n642 ) );
  NOR4_X1 us12_U127 (.A4( us12_n470 ) , .ZN( us12_n476 ) , .A3( us12_n556 ) , .A1( us12_n735 ) , .A2( us12_n755 ) );
  NOR4_X1 us12_U128 (.ZN( us12_n474 ) , .A1( us12_n506 ) , .A3( us12_n544 ) , .A2( us12_n583 ) , .A4( us12_n716 ) );
  NOR2_X1 us12_U129 (.ZN( us12_n733 ) , .A2( us12_n832 ) , .A1( us12_n845 ) );
  NOR2_X1 us12_U13 (.ZN( us12_n495 ) , .A1( us12_n678 ) , .A2( us12_n694 ) );
  NOR2_X1 us12_U130 (.ZN( us12_n789 ) , .A2( us12_n862 ) , .A1( us12_n868 ) );
  NAND4_X1 us12_U131 (.A4( us12_n573 ) , .A3( us12_n574 ) , .A1( us12_n575 ) , .ZN( us12_n723 ) , .A2( us12_n874 ) );
  NOR4_X1 us12_U132 (.A4( us12_n569 ) , .A3( us12_n570 ) , .A2( us12_n571 ) , .A1( us12_n572 ) , .ZN( us12_n573 ) );
  AOI221_X1 us12_U133 (.A( us12_n564 ) , .C2( us12_n565 ) , .ZN( us12_n574 ) , .B2( us12_n845 ) , .B1( us12_n852 ) , .C1( us12_n853 ) );
  NOR2_X1 us12_U134 (.ZN( us12_n575 ) , .A1( us12_n622 ) , .A2( us12_n745 ) );
  NAND4_X1 us12_U135 (.A4( us12_n633 ) , .A3( us12_n634 ) , .A2( us12_n635 ) , .A1( us12_n636 ) , .ZN( us12_n743 ) );
  AOI211_X1 us12_U136 (.B( us12_n623 ) , .A( us12_n624 ) , .ZN( us12_n635 ) , .C2( us12_n836 ) , .C1( us12_n863 ) );
  NOR4_X1 us12_U137 (.A4( us12_n629 ) , .A3( us12_n630 ) , .A2( us12_n631 ) , .A1( us12_n632 ) , .ZN( us12_n633 ) );
  NOR4_X1 us12_U138 (.A4( us12_n626 ) , .A3( us12_n627 ) , .A2( us12_n628 ) , .ZN( us12_n634 ) , .A1( us12_n664 ) );
  NAND4_X1 us12_U139 (.A4( us12_n493 ) , .A3( us12_n494 ) , .A1( us12_n495 ) , .ZN( us12_n802 ) , .A2( us12_n867 ) );
  NOR2_X1 us12_U14 (.A1( us12_n678 ) , .ZN( us12_n693 ) , .A2( us12_n807 ) );
  AOI221_X1 us12_U140 (.A( us12_n489 ) , .ZN( us12_n494 ) , .B2( us12_n836 ) , .C2( us12_n841 ) , .C1( us12_n851 ) , .B1( us12_n860 ) );
  INV_X1 us12_U141 (.A( us12_n778 ) , .ZN( us12_n867 ) );
  NOR4_X1 us12_U142 (.A2( us12_n491 ) , .A1( us12_n492 ) , .ZN( us12_n493 ) , .A3( us12_n580 ) , .A4( us12_n612 ) );
  NOR4_X1 us12_U143 (.A3( us12_n755 ) , .A2( us12_n756 ) , .A1( us12_n757 ) , .ZN( us12_n758 ) , .A4( us12_n869 ) );
  AOI211_X1 us12_U144 (.B( us12_n745 ) , .A( us12_n746 ) , .ZN( us12_n759 ) , .C1( us12_n832 ) , .C2( us12_n853 ) );
  NOR3_X1 us12_U145 (.A3( us12_n741 ) , .A2( us12_n742 ) , .A1( us12_n743 ) , .ZN( us12_n760 ) );
  NOR2_X1 us12_U146 (.ZN( us12_n647 ) , .A1( us12_n854 ) , .A2( us12_n868 ) );
  INV_X1 us12_U147 (.A( us12_n762 ) , .ZN( us12_n830 ) );
  INV_X1 us12_U148 (.A( us12_n754 ) , .ZN( us12_n869 ) );
  OAI21_X1 us12_U149 (.B1( us12_n753 ) , .ZN( us12_n754 ) , .A( us12_n845 ) , .B2( us12_n868 ) );
  INV_X1 us12_U15 (.A( us12_n607 ) , .ZN( us12_n874 ) );
  OR4_X1 us12_U150 (.ZN( us12_n466 ) , .A4( us12_n518 ) , .A3( us12_n529 ) , .A2( us12_n578 ) , .A1( us12_n712 ) );
  OR4_X1 us12_U151 (.A4( us12_n566 ) , .A3( us12_n567 ) , .A2( us12_n568 ) , .ZN( us12_n572 ) , .A1( us12_n665 ) );
  OR4_X1 us12_U152 (.ZN( us12_n492 ) , .A4( us12_n534 ) , .A2( us12_n547 ) , .A1( us12_n559 ) , .A3( us12_n632 ) );
  OR4_X1 us12_U153 (.A4( us12_n518 ) , .A2( us12_n519 ) , .A1( us12_n520 ) , .ZN( us12_n522 ) , .A3( us12_n821 ) );
  OR4_X1 us12_U154 (.A4( us12_n682 ) , .A3( us12_n683 ) , .A2( us12_n684 ) , .A1( us12_n685 ) , .ZN( us12_n690 ) );
  OR4_X1 us12_U155 (.A4( us12_n580 ) , .A3( us12_n581 ) , .A2( us12_n582 ) , .A1( us12_n583 ) , .ZN( us12_n584 ) );
  NAND2_X1 us12_U156 (.ZN( us12_n613 ) , .A2( us12_n837 ) , .A1( us12_n873 ) );
  OR3_X1 us12_U157 (.A3( us12_n506 ) , .A2( us12_n507 ) , .A1( us12_n508 ) , .ZN( us12_n511 ) );
  INV_X1 us12_U158 (.A( us12_n463 ) , .ZN( us12_n864 ) );
  OAI21_X1 us12_U159 (.ZN( us12_n463 ) , .B1( us12_n809 ) , .A( us12_n834 ) , .B2( us12_n851 ) );
  INV_X1 us12_U16 (.A( us12_n680 ) , .ZN( us12_n840 ) );
  INV_X1 us12_U160 (.A( us12_n672 ) , .ZN( us12_n859 ) );
  AOI21_X1 us12_U161 (.A( us12_n670 ) , .B1( us12_n671 ) , .ZN( us12_n672 ) , .B2( us12_n856 ) );
  OAI222_X1 us12_U162 (.B2( us12_n708 ) , .ZN( us12_n709 ) , .C2( us12_n724 ) , .B1( us12_n747 ) , .A1( us12_n806 ) , .C1( us12_n814 ) , .A2( us12_n815 ) );
  AOI22_X1 us12_U163 (.ZN( us12_n696 ) , .A1( us12_n830 ) , .B2( us12_n843 ) , .A2( us12_n865 ) , .B1( us12_n868 ) );
  INV_X1 us12_U164 (.A( us12_n730 ) , .ZN( us12_n839 ) );
  NAND2_X1 us12_U165 (.A1( us12_n447 ) , .A2( us12_n465 ) , .ZN( us12_n749 ) );
  AOI221_X1 us12_U166 (.A( us12_n483 ) , .ZN( us12_n488 ) , .B1( us12_n831 ) , .C2( us12_n844 ) , .C1( us12_n852 ) , .B2( us12_n862 ) );
  OAI22_X1 us12_U167 (.ZN( us12_n483 ) , .A1( us12_n708 ) , .B2( us12_n785 ) , .A2( us12_n806 ) , .B1( us12_n812 ) );
  INV_X1 us12_U168 (.A( us12_n790 ) , .ZN( us12_n832 ) );
  NAND2_X1 us12_U169 (.A1( us12_n451 ) , .A2( us12_n453 ) , .ZN( us12_n762 ) );
  NOR4_X1 us12_U17 (.A4( us12_n445 ) , .A3( us12_n446 ) , .A2( us12_n516 ) , .A1( us12_n541 ) , .ZN( us12_n706 ) );
  AOI211_X1 us12_U170 (.A( us12_n637 ) , .ZN( us12_n645 ) , .B( us12_n743 ) , .C2( us12_n839 ) , .C1( us12_n854 ) );
  OAI22_X1 us12_U171 (.ZN( us12_n637 ) , .A1( us12_n699 ) , .B2( us12_n728 ) , .A2( us12_n762 ) , .B1( us12_n816 ) );
  INV_X1 us12_U172 (.A( us12_n786 ) , .ZN( us12_n862 ) );
  OAI22_X1 us12_U173 (.B2( us12_n779 ) , .B1( us12_n780 ) , .ZN( us12_n781 ) , .A2( us12_n814 ) , .A1( us12_n815 ) );
  OAI22_X1 us12_U174 (.ZN( us12_n489 ) , .A1( us12_n724 ) , .B2( us12_n728 ) , .B1( us12_n730 ) , .A2( us12_n779 ) );
  INV_X1 us12_U175 (.A( us12_n788 ) , .ZN( us12_n845 ) );
  INV_X1 us12_U176 (.A( us12_n816 ) , .ZN( us12_n831 ) );
  OAI22_X1 us12_U177 (.A1( us12_n724 ) , .ZN( us12_n726 ) , .B2( us12_n750 ) , .B1( us12_n812 ) , .A2( us12_n816 ) );
  OAI22_X1 us12_U178 (.B2( us12_n803 ) , .B1( us12_n804 ) , .A2( us12_n805 ) , .A1( us12_n806 ) , .ZN( us12_n808 ) );
  OAI22_X1 us12_U179 (.ZN( us12_n496 ) , .A2( us12_n744 ) , .A1( us12_n780 ) , .B1( us12_n791 ) , .B2( us12_n806 ) );
  OR3_X1 us12_U18 (.ZN( us12_n446 ) , .A1( us12_n528 ) , .A3( us12_n577 ) , .A2( us12_n875 ) );
  INV_X1 us12_U180 (.A( us12_n814 ) , .ZN( us12_n833 ) );
  INV_X1 us12_U181 (.A( us12_n805 ) , .ZN( us12_n860 ) );
  OAI22_X1 us12_U182 (.ZN( us12_n710 ) , .A2( us12_n728 ) , .B2( us12_n729 ) , .A1( us12_n744 ) , .B1( us12_n813 ) );
  INV_X1 us12_U183 (.A( us12_n750 ) , .ZN( us12_n842 ) );
  OAI22_X1 us12_U184 (.B1( us12_n490 ) , .ZN( us12_n491 ) , .A1( us12_n686 ) , .A2( us12_n763 ) , .B2( us12_n817 ) );
  NOR3_X1 us12_U185 (.ZN( us12_n490 ) , .A1( us12_n782 ) , .A2( us12_n850 ) , .A3( us12_n863 ) );
  OAI22_X1 us12_U186 (.ZN( us12_n695 ) , .A2( us12_n730 ) , .A1( us12_n780 ) , .B1( us12_n791 ) , .B2( us12_n817 ) );
  OAI22_X1 us12_U187 (.B2( us12_n744 ) , .ZN( us12_n746 ) , .A2( us12_n762 ) , .B1( us12_n780 ) , .A1( us12_n792 ) );
  NOR2_X1 us12_U188 (.ZN( us12_n532 ) , .A2( us12_n749 ) , .A1( us12_n750 ) );
  INV_X1 us12_U189 (.A( us12_n744 ) , .ZN( us12_n837 ) );
  OR4_X1 us12_U19 (.A4( us12_n442 ) , .A2( us12_n443 ) , .A1( us12_n444 ) , .ZN( us12_n445 ) , .A3( us12_n553 ) );
  NOR2_X1 us12_U190 (.ZN( us12_n666 ) , .A1( us12_n728 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U191 (.ZN( us12_n615 ) , .A1( us12_n785 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U192 (.ZN( us12_n629 ) , .A2( us12_n728 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U193 (.ZN( us12_n715 ) , .A1( us12_n805 ) , .A2( us12_n817 ) );
  NOR2_X1 us12_U194 (.ZN( us12_n570 ) , .A1( us12_n728 ) , .A2( us12_n806 ) );
  NOR2_X1 us12_U195 (.A2( us12_n708 ) , .A1( us12_n750 ) , .ZN( us12_n771 ) );
  NOR2_X1 us12_U196 (.ZN( us12_n611 ) , .A2( us12_n780 ) , .A1( us12_n806 ) );
  NOR2_X1 us12_U197 (.ZN( us12_n601 ) , .A2( us12_n780 ) , .A1( us12_n803 ) );
  NOR2_X1 us12_U198 (.ZN( us12_n667 ) , .A1( us12_n750 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U199 (.ZN( us12_n555 ) , .A1( us12_n750 ) , .A2( us12_n791 ) );
  INV_X1 us12_U20 (.A( us12_n613 ) , .ZN( us12_n875 ) );
  NOR2_X1 us12_U200 (.ZN( us12_n654 ) , .A1( us12_n728 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U201 (.ZN( us12_n528 ) , .A2( us12_n724 ) , .A1( us12_n803 ) );
  NOR2_X1 us12_U202 (.ZN( us12_n546 ) , .A2( us12_n780 ) , .A1( us12_n814 ) );
  NOR2_X1 us12_U203 (.ZN( us12_n577 ) , .A2( us12_n699 ) , .A1( us12_n814 ) );
  NOR2_X1 us12_U204 (.ZN( us12_n508 ) , .A2( us12_n780 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U205 (.ZN( us12_n543 ) , .A2( us12_n708 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U206 (.ZN( us12_n664 ) , .A1( us12_n785 ) , .A2( us12_n791 ) );
  NOR2_X1 us12_U207 (.A2( us12_n744 ) , .ZN( us12_n755 ) , .A1( us12_n805 ) );
  NOR2_X1 us12_U208 (.ZN( us12_n735 ) , .A2( us12_n803 ) , .A1( us12_n805 ) );
  INV_X1 us12_U209 (.A( us12_n792 ) , .ZN( us12_n851 ) );
  INV_X1 us12_U21 (.A( us12_n749 ) , .ZN( us12_n863 ) );
  INV_X1 us12_U210 (.A( us12_n728 ) , .ZN( us12_n852 ) );
  NOR2_X1 us12_U211 (.A2( us12_n744 ) , .ZN( us12_n769 ) , .A1( us12_n812 ) );
  INV_X1 us12_U212 (.A( us12_n747 ) , .ZN( us12_n834 ) );
  NOR2_X1 us12_U213 (.A1( us12_n699 ) , .ZN( us12_n768 ) , .A2( us12_n813 ) );
  INV_X1 us12_U214 (.A( us12_n806 ) , .ZN( us12_n841 ) );
  NOR2_X1 us12_U215 (.ZN( us12_n531 ) , .A2( us12_n780 ) , .A1( us12_n816 ) );
  NOR2_X1 us12_U216 (.ZN( us12_n509 ) , .A1( us12_n729 ) , .A2( us12_n779 ) );
  NOR2_X1 us12_U217 (.ZN( us12_n599 ) , .A2( us12_n791 ) , .A1( us12_n816 ) );
  NOR2_X1 us12_U218 (.ZN( us12_n661 ) , .A1( us12_n729 ) , .A2( us12_n790 ) );
  NOR2_X1 us12_U219 (.ZN( us12_n507 ) , .A1( us12_n812 ) , .A2( us12_n817 ) );
  AOI222_X1 us12_U22 (.ZN( us12_n605 ) , .B2( us12_n671 ) , .B1( us12_n753 ) , .C2( us12_n831 ) , .A1( us12_n833 ) , .A2( us12_n862 ) , .C1( us12_n863 ) );
  NOR2_X1 us12_U220 (.ZN( us12_n544 ) , .A2( us12_n785 ) , .A1( us12_n792 ) );
  NOR2_X1 us12_U221 (.A1( us12_n749 ) , .ZN( us12_n767 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U222 (.ZN( us12_n545 ) , .A1( us12_n749 ) , .A2( us12_n814 ) );
  NOR2_X1 us12_U223 (.ZN( us12_n557 ) , .A1( us12_n792 ) , .A2( us12_n814 ) );
  NOR2_X1 us12_U224 (.ZN( us12_n556 ) , .A1( us12_n762 ) , .A2( us12_n805 ) );
  NOR2_X1 us12_U225 (.ZN( us12_n609 ) , .A2( us12_n724 ) , .A1( us12_n817 ) );
  NOR2_X1 us12_U226 (.ZN( us12_n663 ) , .A1( us12_n729 ) , .A2( us12_n785 ) );
  NOR2_X1 us12_U227 (.ZN( us12_n517 ) , .A1( us12_n708 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U228 (.ZN( us12_n506 ) , .A2( us12_n728 ) , .A1( us12_n762 ) );
  OAI22_X1 us12_U229 (.B1( us12_n440 ) , .ZN( us12_n444 ) , .A2( us12_n728 ) , .A1( us12_n744 ) , .B2( us12_n749 ) );
  AOI222_X1 us12_U23 (.ZN( us12_n563 ) , .B1( us12_n830 ) , .C1( us12_n841 ) , .A2( us12_n843 ) , .A1( us12_n854 ) , .B2( us12_n863 ) , .C2( us12_n873 ) );
  NOR3_X1 us12_U230 (.ZN( us12_n440 ) , .A2( us12_n836 ) , .A3( us12_n837 ) , .A1( us12_n846 ) );
  NOR2_X1 us12_U231 (.ZN( us12_n614 ) , .A1( us12_n762 ) , .A2( us12_n812 ) );
  NOR2_X1 us12_U232 (.ZN( us12_n533 ) , .A2( us12_n724 ) , .A1( us12_n730 ) );
  NOR2_X1 us12_U233 (.ZN( us12_n579 ) , .A2( us12_n708 ) , .A1( us12_n730 ) );
  NOR2_X1 us12_U234 (.ZN( us12_n521 ) , .A1( us12_n790 ) , .A2( us12_n812 ) );
  NOR2_X1 us12_U235 (.ZN( us12_n558 ) , .A1( us12_n708 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U236 (.ZN( us12_n655 ) , .A1( us12_n790 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U237 (.ZN( us12_n670 ) , .A1( us12_n790 ) , .A2( us12_n805 ) );
  NOR2_X1 us12_U238 (.ZN( us12_n668 ) , .A2( us12_n708 ) , .A1( us12_n790 ) );
  NOR2_X1 us12_U239 (.ZN( us12_n530 ) , .A2( us12_n744 ) , .A1( us12_n792 ) );
  AOI222_X1 us12_U24 (.ZN( us12_n660 ) , .A2( us12_n839 ) , .B1( us12_n841 ) , .C2( us12_n845 ) , .A1( us12_n860 ) , .C1( us12_n863 ) , .B2( us12_n870 ) );
  NOR2_X1 us12_U240 (.ZN( us12_n631 ) , .A1( us12_n724 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U241 (.ZN( us12_n630 ) , .A1( us12_n747 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U242 (.ZN( us12_n542 ) , .A1( us12_n762 ) , .A2( us12_n791 ) );
  INV_X1 us12_U243 (.A( us12_n763 ) , .ZN( us12_n866 ) );
  AOI21_X1 us12_U244 (.ZN( us12_n515 ) , .A( us12_n729 ) , .B1( us12_n750 ) , .B2( us12_n803 ) );
  NOR2_X1 us12_U245 (.ZN( us12_n718 ) , .A2( us12_n724 ) , .A1( us12_n744 ) );
  NOR2_X1 us12_U246 (.ZN( us12_n516 ) , .A1( us12_n708 ) , .A2( us12_n744 ) );
  INV_X1 us12_U247 (.A( us12_n729 ) , .ZN( us12_n868 ) );
  NOR2_X1 us12_U248 (.ZN( us12_n656 ) , .A1( us12_n747 ) , .A2( us12_n780 ) );
  AOI21_X1 us12_U249 (.ZN( us12_n540 ) , .A( us12_n763 ) , .B2( us12_n779 ) , .B1( us12_n817 ) );
  INV_X1 us12_U25 (.A( us12_n647 ) , .ZN( us12_n870 ) );
  NOR2_X1 us12_U250 (.ZN( us12_n559 ) , .A2( us12_n791 ) , .A1( us12_n803 ) );
  NOR2_X1 us12_U251 (.A2( us12_n708 ) , .A1( us12_n762 ) , .ZN( us12_n794 ) );
  NOR2_X1 us12_U252 (.ZN( us12_n642 ) , .A2( us12_n788 ) , .A1( us12_n791 ) );
  NOR2_X1 us12_U253 (.ZN( us12_n683 ) , .A2( us12_n699 ) , .A1( us12_n803 ) );
  AOI21_X1 us12_U254 (.B1( us12_n625 ) , .ZN( us12_n627 ) , .A( us12_n763 ) , .B2( us12_n814 ) );
  AOI21_X1 us12_U255 (.A( us12_n815 ) , .B2( us12_n816 ) , .B1( us12_n817 ) , .ZN( us12_n818 ) );
  AOI21_X1 us12_U256 (.ZN( us12_n650 ) , .A( us12_n779 ) , .B1( us12_n792 ) , .B2( us12_n805 ) );
  AOI21_X1 us12_U257 (.ZN( us12_n499 ) , .B1( us12_n680 ) , .A( us12_n812 ) , .B2( us12_n816 ) );
  NOR2_X1 us12_U258 (.ZN( us12_n520 ) , .A2( us12_n708 ) , .A1( us12_n814 ) );
  AOI21_X1 us12_U259 (.ZN( us12_n569 ) , .B1( us12_n750 ) , .B2( us12_n762 ) , .A( us12_n780 ) );
  NOR4_X1 us12_U26 (.ZN( us12_n473 ) , .A2( us12_n521 ) , .A4( us12_n594 ) , .A1( us12_n609 ) , .A3( us12_n629 ) );
  OAI221_X1 us12_U260 (.A( us12_n727 ) , .C2( us12_n728 ) , .B2( us12_n729 ) , .B1( us12_n730 ) , .ZN( us12_n737 ) , .C1( us12_n817 ) );
  AOI22_X1 us12_U261 (.ZN( us12_n727 ) , .B1( us12_n832 ) , .A2( us12_n838 ) , .A1( us12_n863 ) , .B2( us12_n866 ) );
  AOI21_X1 us12_U262 (.ZN( us12_n589 ) , .B2( us12_n699 ) , .B1( us12_n815 ) , .A( us12_n817 ) );
  NOR2_X1 us12_U263 (.ZN( us12_n519 ) , .A2( us12_n699 ) , .A1( us12_n816 ) );
  AOI21_X1 us12_U264 (.ZN( us12_n539 ) , .B2( us12_n812 ) , .A( us12_n814 ) , .B1( us12_n815 ) );
  AOI21_X1 us12_U265 (.ZN( us12_n640 ) , .B2( us12_n747 ) , .A( us12_n792 ) , .B1( us12_n803 ) );
  AOI21_X1 us12_U266 (.ZN( us12_n514 ) , .A( us12_n779 ) , .B2( us12_n792 ) , .B1( us12_n812 ) );
  AOI21_X1 us12_U267 (.B1( us12_n699 ) , .ZN( us12_n700 ) , .A( us12_n732 ) , .B2( us12_n763 ) );
  AOI21_X1 us12_U268 (.ZN( us12_n591 ) , .B2( us12_n763 ) , .A( us12_n785 ) , .B1( us12_n812 ) );
  AOI21_X1 us12_U269 (.ZN( us12_n593 ) , .B1( us12_n750 ) , .A( us12_n792 ) , .B2( us12_n813 ) );
  NOR4_X1 us12_U27 (.A4( us12_n544 ) , .A3( us12_n545 ) , .A2( us12_n546 ) , .A1( us12_n547 ) , .ZN( us12_n548 ) );
  NOR2_X1 us12_U270 (.ZN( us12_n547 ) , .A1( us12_n699 ) , .A2( us12_n744 ) );
  INV_X1 us12_U271 (.A( us12_n791 ) , .ZN( us12_n873 ) );
  AOI21_X1 us12_U272 (.ZN( us12_n564 ) , .B1( us12_n724 ) , .A( us12_n779 ) , .B2( us12_n791 ) );
  AOI21_X1 us12_U273 (.ZN( us12_n497 ) , .A( us12_n779 ) , .B2( us12_n791 ) , .B1( us12_n804 ) );
  AOI21_X1 us12_U274 (.ZN( us12_n498 ) , .A( us12_n724 ) , .B2( us12_n762 ) , .B1( us12_n814 ) );
  AOI21_X1 us12_U275 (.ZN( us12_n649 ) , .B1( us12_n729 ) , .B2( us12_n763 ) , .A( us12_n813 ) );
  NOR2_X1 us12_U276 (.ZN( us12_n529 ) , .A1( us12_n708 ) , .A2( us12_n779 ) );
  NOR2_X1 us12_U277 (.ZN( us12_n685 ) , .A1( us12_n729 ) , .A2( us12_n816 ) );
  AOI21_X1 us12_U278 (.B1( us12_n686 ) , .ZN( us12_n687 ) , .A( us12_n728 ) , .B2( us12_n761 ) );
  AOI21_X1 us12_U279 (.A( us12_n812 ) , .B2( us12_n813 ) , .B1( us12_n814 ) , .ZN( us12_n819 ) );
  NOR4_X1 us12_U28 (.A4( us12_n532 ) , .A3( us12_n533 ) , .A2( us12_n534 ) , .ZN( us12_n535 ) , .A1( us12_n820 ) );
  AOI21_X1 us12_U280 (.ZN( us12_n450 ) , .B2( us12_n792 ) , .A( us12_n803 ) , .B1( us12_n815 ) );
  NOR2_X1 us12_U281 (.ZN( us12_n568 ) , .A1( us12_n729 ) , .A2( us12_n762 ) );
  NOR2_X1 us12_U282 (.ZN( us12_n682 ) , .A2( us12_n708 ) , .A1( us12_n817 ) );
  AOI21_X1 us12_U283 (.ZN( us12_n641 ) , .B1( us12_n680 ) , .A( us12_n791 ) , .B2( us12_n817 ) );
  INV_X1 us12_U284 (.A( us12_n699 ) , .ZN( us12_n853 ) );
  AOI21_X1 us12_U285 (.ZN( us12_n689 ) , .B2( us12_n749 ) , .B1( us12_n763 ) , .A( us12_n806 ) );
  AOI21_X1 us12_U286 (.ZN( us12_n639 ) , .B2( us12_n749 ) , .A( us12_n788 ) , .B1( us12_n812 ) );
  AOI21_X1 us12_U287 (.A( us12_n790 ) , .B2( us12_n791 ) , .B1( us12_n792 ) , .ZN( us12_n793 ) );
  AOI21_X1 us12_U288 (.A( us12_n733 ) , .ZN( us12_n734 ) , .B2( us12_n780 ) , .B1( us12_n792 ) );
  NOR2_X1 us12_U289 (.ZN( us12_n567 ) , .A1( us12_n747 ) , .A2( us12_n805 ) );
  NOR4_X1 us12_U29 (.ZN( us12_n479 ) , .A1( us12_n520 ) , .A4( us12_n557 ) , .A3( us12_n582 ) , .A2( us12_n630 ) );
  NAND2_X1 us12_U290 (.ZN( us12_n753 ) , .A1( us12_n763 ) , .A2( us12_n805 ) );
  NOR2_X1 us12_U291 (.A2( us12_n813 ) , .A1( us12_n815 ) , .ZN( us12_n821 ) );
  NOR2_X1 us12_U292 (.ZN( us12_n578 ) , .A1( us12_n708 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U293 (.ZN( us12_n665 ) , .A1( us12_n780 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U294 (.ZN( us12_n711 ) , .A1( us12_n762 ) , .A2( us12_n763 ) );
  NOR2_X1 us12_U295 (.ZN( us12_n583 ) , .A1( us12_n792 ) , .A2( us12_n817 ) );
  AOI21_X1 us12_U296 (.ZN( us12_n442 ) , .A( us12_n699 ) , .B1( us12_n733 ) , .B2( us12_n750 ) );
  NOR2_X1 us12_U297 (.ZN( us12_n534 ) , .A1( us12_n724 ) , .A2( us12_n788 ) );
  NOR2_X1 us12_U298 (.ZN( us12_n582 ) , .A1( us12_n744 ) , .A2( us12_n815 ) );
  NOR2_X1 us12_U299 (.ZN( us12_n684 ) , .A1( us12_n791 ) , .A2( us12_n813 ) );
  NAND2_X1 us12_U3 (.A1( us12_n449 ) , .A2( us12_n460 ) , .ZN( us12_n792 ) );
  NOR4_X1 us12_U30 (.ZN( us12_n456 ) , .A2( us12_n517 ) , .A1( us12_n543 ) , .A3( us12_n579 ) , .A4( us12_n615 ) );
  OAI21_X1 us12_U300 (.A( us12_n698 ) , .ZN( us12_n702 ) , .B2( us12_n750 ) , .B1( us12_n804 ) );
  OAI21_X1 us12_U301 (.ZN( us12_n698 ) , .B2( us12_n833 ) , .B1( us12_n838 ) , .A( us12_n860 ) );
  INV_X1 us12_U302 (.A( us12_n815 ) , .ZN( us12_n855 ) );
  INV_X1 us12_U303 (.A( us12_n785 ) , .ZN( us12_n846 ) );
  OAI21_X1 us12_U304 (.A( us12_n731 ) , .B1( us12_n732 ) , .ZN( us12_n736 ) , .B2( us12_n805 ) );
  OAI21_X1 us12_U305 (.ZN( us12_n731 ) , .A( us12_n833 ) , .B2( us12_n852 ) , .B1( us12_n873 ) );
  INV_X1 us12_U306 (.A( us12_n780 ) , .ZN( us12_n850 ) );
  INV_X1 us12_U307 (.A( us12_n813 ) , .ZN( us12_n836 ) );
  OAI221_X1 us12_U308 (.A( us12_n783 ) , .C2( us12_n784 ) , .B2( us12_n785 ) , .B1( us12_n786 ) , .ZN( us12_n796 ) , .C1( us12_n813 ) );
  AOI22_X1 us12_U309 (.A2( us12_n782 ) , .ZN( us12_n783 ) , .B2( us12_n831 ) , .A1( us12_n834 ) , .B1( us12_n863 ) );
  AOI221_X1 us12_U31 (.A( us12_n713 ) , .B2( us12_n714 ) , .ZN( us12_n720 ) , .C1( us12_n832 ) , .B1( us12_n839 ) , .C2( us12_n863 ) );
  OAI21_X1 us12_U310 (.A( us12_n787 ) , .B2( us12_n788 ) , .B1( us12_n789 ) , .ZN( us12_n795 ) );
  OAI21_X1 us12_U311 (.ZN( us12_n787 ) , .A( us12_n839 ) , .B1( us12_n863 ) , .B2( us12_n873 ) );
  NAND2_X1 us12_U312 (.A2( us12_n762 ) , .A1( us12_n806 ) , .ZN( us12_n810 ) );
  NOR2_X1 us12_U313 (.ZN( us12_n470 ) , .A2( us12_n779 ) , .A1( us12_n815 ) );
  NOR2_X1 us12_U314 (.ZN( us12_n484 ) , .A1( us12_n788 ) , .A2( us12_n805 ) );
  NAND2_X1 us12_U315 (.ZN( us12_n714 ) , .A1( us12_n728 ) , .A2( us12_n780 ) );
  NAND2_X1 us12_U316 (.ZN( us12_n671 ) , .A1( us12_n806 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U317 (.ZN( us12_n526 ) , .A1( us12_n724 ) , .A2( us12_n750 ) );
  AOI21_X1 us12_U318 (.ZN( us12_n443 ) , .B1( us12_n789 ) , .B2( us12_n791 ) , .A( us12_n814 ) );
  INV_X1 us12_U319 (.A( us12_n817 ) , .ZN( us12_n844 ) );
  OR2_X1 us12_U32 (.A2( us12_n711 ) , .A1( us12_n712 ) , .ZN( us12_n713 ) );
  NOR2_X1 us12_U320 (.ZN( us12_n712 ) , .A2( us12_n724 ) , .A1( us12_n790 ) );
  NAND2_X1 us12_U321 (.A1( us12_n699 ) , .A2( us12_n729 ) , .ZN( us12_n782 ) );
  NOR2_X1 us12_U322 (.ZN( us12_n518 ) , .A1( us12_n708 ) , .A2( us12_n788 ) );
  OAI22_X1 us12_U323 (.B2( us12_n750 ) , .B1( us12_n751 ) , .A1( us12_n752 ) , .ZN( us12_n756 ) , .A2( us12_n806 ) );
  NOR3_X1 us12_U324 (.ZN( us12_n752 ) , .A2( us12_n853 ) , .A1( us12_n863 ) , .A3( us12_n865 ) );
  NOR2_X1 us12_U325 (.ZN( us12_n751 ) , .A2( us12_n852 ) , .A1( us12_n860 ) );
  INV_X1 us12_U326 (.A( us12_n724 ) , .ZN( us12_n856 ) );
  NAND2_X2 us12_U327 (.A2( us12_n454 ) , .A1( us12_n472 ) , .ZN( us12_n779 ) );
  AND2_X1 us12_U328 (.ZN( us12_n732 ) , .A1( us12_n779 ) , .A2( us12_n785 ) );
  AOI221_X1 us12_U329 (.A( us12_n764 ) , .ZN( us12_n774 ) , .C2( us12_n810 ) , .B2( us12_n835 ) , .C1( us12_n855 ) , .B1( us12_n866 ) );
  NOR2_X1 us12_U33 (.ZN( us12_n680 ) , .A2( us12_n834 ) , .A1( us12_n839 ) );
  AOI21_X1 us12_U330 (.B2( us12_n763 ) , .ZN( us12_n764 ) , .A( us12_n788 ) , .B1( us12_n792 ) );
  INV_X1 us12_U331 (.A( us12_n761 ) , .ZN( us12_n835 ) );
  NAND2_X1 us12_U332 (.A2( us12_n448 ) , .A1( us12_n460 ) , .ZN( us12_n728 ) );
  NAND2_X1 us12_U333 (.A1( us12_n451 ) , .A2( us12_n454 ) , .ZN( us12_n814 ) );
  NAND2_X1 us12_U334 (.A1( us12_n447 ) , .A2( us12_n449 ) , .ZN( us12_n805 ) );
  NAND2_X1 us12_U335 (.A1( us12_n451 ) , .A2( us12_n471 ) , .ZN( us12_n816 ) );
  NAND2_X1 us12_U336 (.A2( us12_n453 ) , .A1( us12_n455 ) , .ZN( us12_n806 ) );
  NAND2_X1 us12_U337 (.A2( us12_n464 ) , .A1( us12_n465 ) , .ZN( us12_n812 ) );
  NAND2_X1 us12_U338 (.A1( us12_n441 ) , .A2( us12_n460 ) , .ZN( us12_n699 ) );
  NAND2_X1 us12_U339 (.A2( us12_n449 ) , .A1( us12_n452 ) , .ZN( us12_n763 ) );
  AOI222_X1 us12_U34 (.ZN( us12_n469 ) , .B1( us12_n832 ) , .A1( us12_n839 ) , .C1( us12_n842 ) , .C2( us12_n851 ) , .A2( us12_n855 ) , .B2( us12_n865 ) );
  NAND2_X2 us12_U340 (.A1( us12_n455 ) , .A2( us12_n462 ) , .ZN( us12_n750 ) );
  NAND2_X1 us12_U341 (.A2( us12_n448 ) , .A1( us12_n452 ) , .ZN( us12_n729 ) );
  NOR2_X1 us12_U342 (.ZN( us12_n453 ) , .A1( us12_n826 ) , .A2( us12_n827 ) );
  NOR2_X1 us12_U343 (.ZN( us12_n465 ) , .A2( us12_n847 ) , .A1( us12_n848 ) );
  NOR2_X1 us12_U344 (.ZN( us12_n451 ) , .A1( us12_n828 ) , .A2( us12_n829 ) );
  NAND2_X1 us12_U345 (.A1( us12_n462 ) , .A2( us12_n472 ) , .ZN( us12_n788 ) );
  NAND2_X1 us12_U346 (.A2( us12_n461 ) , .A1( us12_n471 ) , .ZN( us12_n697 ) );
  NAND2_X1 us12_U347 (.A2( us12_n461 ) , .A1( us12_n462 ) , .ZN( us12_n747 ) );
  NAND2_X1 us12_U348 (.A1( us12_n451 ) , .A2( us12_n462 ) , .ZN( us12_n790 ) );
  NAND2_X1 us12_U349 (.A1( us12_n452 ) , .A2( us12_n465 ) , .ZN( us12_n669 ) );
  NOR4_X1 us12_U35 (.A1( us12_n466 ) , .ZN( us12_n467 ) , .A4( us12_n542 ) , .A2( us12_n554 ) , .A3( us12_n614 ) );
  NAND2_X1 us12_U350 (.A2( us12_n441 ) , .A1( us12_n447 ) , .ZN( us12_n784 ) );
  NAND2_X2 us12_U351 (.A1( us12_n441 ) , .A2( us12_n464 ) , .ZN( us12_n708 ) );
  NAND2_X1 us12_U352 (.A2( us12_n471 ) , .A1( us12_n472 ) , .ZN( us12_n817 ) );
  NAND2_X1 us12_U353 (.A2( us12_n454 ) , .A1( us12_n455 ) , .ZN( us12_n730 ) );
  NOR2_X1 us12_U354 (.ZN( us12_n447 ) , .A2( us12_n849 ) , .A1( us12_n858 ) );
  NAND2_X1 us12_U355 (.A1( us12_n447 ) , .A2( us12_n448 ) , .ZN( us12_n786 ) );
  NAND2_X1 us12_U356 (.A1( us12_n454 ) , .A2( us12_n461 ) , .ZN( us12_n813 ) );
  NAND2_X2 us12_U357 (.A1( us12_n453 ) , .A2( us12_n472 ) , .ZN( us12_n785 ) );
  NAND2_X1 us12_U358 (.A1( us12_n453 ) , .A2( us12_n461 ) , .ZN( us12_n744 ) );
  NOR2_X1 us12_U359 (.A2( sa12_6 ) , .A1( sa12_7 ) , .ZN( us12_n464 ) );
  AOI221_X1 us12_U36 (.ZN( us12_n468 ) , .C2( us12_n714 ) , .B2( us12_n831 ) , .C1( us12_n845 ) , .B1( us12_n860 ) , .A( us12_n864 ) );
  NOR2_X1 us12_U360 (.A2( sa12_2 ) , .ZN( us12_n461 ) , .A1( us12_n829 ) );
  NOR2_X1 us12_U361 (.A2( sa12_7 ) , .ZN( us12_n460 ) , .A1( us12_n849 ) );
  NOR2_X1 us12_U362 (.A2( sa12_4 ) , .ZN( us12_n449 ) , .A1( us12_n848 ) );
  NOR2_X1 us12_U363 (.A2( sa12_4 ) , .A1( sa12_5 ) , .ZN( us12_n441 ) );
  NOR2_X1 us12_U364 (.A2( sa12_5 ) , .ZN( us12_n448 ) , .A1( us12_n847 ) );
  NOR2_X1 us12_U365 (.A2( sa12_0 ) , .ZN( us12_n454 ) , .A1( us12_n827 ) );
  NOR2_X1 us12_U366 (.A2( sa12_1 ) , .ZN( us12_n471 ) , .A1( us12_n826 ) );
  NOR2_X1 us12_U367 (.A2( sa12_6 ) , .ZN( us12_n452 ) , .A1( us12_n858 ) );
  NOR2_X1 us12_U368 (.A2( sa12_0 ) , .A1( sa12_1 ) , .ZN( us12_n462 ) );
  INV_X1 us12_U369 (.A( sa12_6 ) , .ZN( us12_n849 ) );
  NOR4_X1 us12_U37 (.A4( us12_n577 ) , .A3( us12_n578 ) , .A2( us12_n579 ) , .ZN( us12_n586 ) , .A1( us12_n683 ) );
  INV_X1 us12_U370 (.A( sa12_4 ) , .ZN( us12_n847 ) );
  INV_X1 us12_U371 (.A( sa12_1 ) , .ZN( us12_n827 ) );
  NAND2_X2 us12_U372 (.A1( us12_n455 ) , .A2( us12_n471 ) , .ZN( us12_n803 ) );
  INV_X1 us12_U373 (.A( sa12_0 ) , .ZN( us12_n826 ) );
  INV_X1 us12_U374 (.A( sa12_7 ) , .ZN( us12_n858 ) );
  INV_X1 us12_U375 (.A( sa12_5 ) , .ZN( us12_n848 ) );
  INV_X1 us12_U376 (.A( sa12_2 ) , .ZN( us12_n828 ) );
  AOI21_X1 us12_U377 (.ZN( us12_n510 ) , .B2( us12_n669 ) , .A( us12_n730 ) , .B1( us12_n815 ) );
  OAI22_X1 us12_U378 (.ZN( us12_n624 ) , .B1( us12_n669 ) , .B2( us12_n747 ) , .A1( us12_n815 ) , .A2( us12_n816 ) );
  AOI21_X1 us12_U379 (.ZN( us12_n626 ) , .B2( us12_n669 ) , .A( us12_n790 ) , .B1( us12_n791 ) );
  NOR4_X1 us12_U38 (.A1( us12_n584 ) , .ZN( us12_n585 ) , .A3( us12_n652 ) , .A2( us12_n662 ) , .A4( us12_n767 ) );
  INV_X1 us12_U380 (.A( us12_n669 ) , .ZN( us12_n865 ) );
  NOR2_X1 us12_U381 (.A1( us12_n669 ) , .ZN( us12_n766 ) , .A2( us12_n813 ) );
  AOI21_X1 us12_U382 (.ZN( us12_n477 ) , .A( us12_n669 ) , .B1( us12_n750 ) , .B2( us12_n806 ) );
  NOR2_X1 us12_U383 (.A1( us12_n669 ) , .ZN( us12_n673 ) , .A2( us12_n744 ) );
  NOR2_X1 us12_U384 (.ZN( us12_n602 ) , .A1( us12_n669 ) , .A2( us12_n803 ) );
  NOR2_X1 us12_U385 (.A1( us12_n669 ) , .ZN( us12_n688 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U386 (.ZN( us12_n527 ) , .A1( us12_n669 ) , .A2( us12_n779 ) );
  NOR2_X1 us12_U387 (.ZN( us12_n652 ) , .A1( us12_n669 ) , .A2( us12_n814 ) );
  NOR2_X1 us12_U388 (.ZN( us12_n628 ) , .A2( us12_n669 ) , .A1( us12_n785 ) );
  NOR2_X1 us12_U389 (.ZN( us12_n581 ) , .A1( us12_n669 ) , .A2( us12_n788 ) );
  NOR4_X1 us12_U39 (.A4( us12_n661 ) , .A3( us12_n662 ) , .A2( us12_n663 ) , .A1( us12_n664 ) , .ZN( us12_n677 ) );
  OAI22_X1 us12_U390 (.ZN( us12_n590 ) , .B1( us12_n730 ) , .B2( us12_n749 ) , .A2( us12_n786 ) , .A1( us12_n803 ) );
  NAND2_X1 us12_U391 (.A2( us12_n749 ) , .A1( us12_n786 ) , .ZN( us12_n809 ) );
  NOR2_X1 us12_U392 (.ZN( us12_n612 ) , .A1( us12_n779 ) , .A2( us12_n786 ) );
  NOR2_X1 us12_U393 (.ZN( us12_n717 ) , .A2( us12_n744 ) , .A1( us12_n786 ) );
  NOR2_X1 us12_U394 (.ZN( us12_n653 ) , .A1( us12_n762 ) , .A2( us12_n786 ) );
  NOR2_X1 us12_U395 (.ZN( us12_n554 ) , .A1( us12_n786 ) , .A2( us12_n813 ) );
  NOR2_X1 us12_U396 (.ZN( us12_n701 ) , .A2( us12_n786 ) , .A1( us12_n817 ) );
  OAI222_X1 us12_U397 (.ZN( us12_n617 ) , .B1( us12_n697 ) , .C1( us12_n724 ) , .C2( us12_n747 ) , .B2( us12_n786 ) , .A2( us12_n792 ) , .A1( us12_n816 ) );
  NOR2_X1 us12_U398 (.A1( us12_n730 ) , .ZN( us12_n765 ) , .A2( us12_n786 ) );
  NAND2_X1 us12_U399 (.A1( us12_n729 ) , .A2( us12_n784 ) , .ZN( us12_n811 ) );
  NAND2_X1 us12_U4 (.A1( us12_n449 ) , .A2( us12_n464 ) , .ZN( us12_n724 ) );
  NOR4_X1 us12_U40 (.A4( us12_n665 ) , .A3( us12_n666 ) , .A2( us12_n667 ) , .A1( us12_n668 ) , .ZN( us12_n676 ) );
  OAI22_X1 us12_U400 (.ZN( us12_n588 ) , .A2( us12_n747 ) , .B2( us12_n762 ) , .A1( us12_n763 ) , .B1( us12_n784 ) );
  OAI221_X1 us12_U401 (.A( us12_n696 ) , .ZN( us12_n703 ) , .C2( us12_n784 ) , .C1( us12_n785 ) , .B1( us12_n786 ) , .B2( us12_n806 ) );
  AOI21_X1 us12_U402 (.ZN( us12_n592 ) , .B1( us12_n728 ) , .B2( us12_n784 ) , .A( us12_n790 ) );
  AOI21_X1 us12_U403 (.ZN( us12_n648 ) , .A( us12_n762 ) , .B2( us12_n784 ) , .B1( us12_n792 ) );
  AOI21_X1 us12_U404 (.ZN( us12_n623 ) , .B1( us12_n699 ) , .A( us12_n779 ) , .B2( us12_n784 ) );
  OAI22_X1 us12_U405 (.ZN( us12_n681 ) , .A1( us12_n699 ) , .A2( us12_n730 ) , .B2( us12_n784 ) , .B1( us12_n817 ) );
  OAI21_X1 us12_U406 (.A( us12_n613 ) , .ZN( us12_n616 ) , .B1( us12_n625 ) , .B2( us12_n784 ) );
  NOR2_X1 us12_U407 (.ZN( us12_n610 ) , .A1( us12_n784 ) , .A2( us12_n816 ) );
  NOR2_X1 us12_U408 (.ZN( us12_n651 ) , .A1( us12_n784 ) , .A2( us12_n788 ) );
  OAI222_X1 us12_U409 (.A2( us12_n669 ) , .ZN( us12_n674 ) , .B1( us12_n747 ) , .B2( us12_n784 ) , .C2( us12_n788 ) , .C1( us12_n815 ) , .A1( us12_n817 ) );
  NOR4_X1 us12_U41 (.A3( us12_n673 ) , .A1( us12_n674 ) , .ZN( us12_n675 ) , .A4( us12_n715 ) , .A2( us12_n859 ) );
  NOR2_X1 us12_U410 (.ZN( us12_n553 ) , .A2( us12_n744 ) , .A1( us12_n784 ) );
  INV_X1 us12_U411 (.A( us12_n784 ) , .ZN( us12_n861 ) );
  AOI21_X1 us12_U412 (.ZN( us12_n500 ) , .A( us12_n697 ) , .B1( us12_n708 ) , .B2( us12_n786 ) );
  INV_X1 us12_U413 (.A( us12_n697 ) , .ZN( us12_n838 ) );
  NOR2_X1 us12_U414 (.A1( us12_n697 ) , .ZN( us12_n770 ) , .A2( us12_n815 ) );
  AOI21_X1 us12_U415 (.ZN( us12_n571 ) , .B2( us12_n697 ) , .B1( us12_n806 ) , .A( us12_n812 ) );
  NOR2_X1 us12_U416 (.ZN( us12_n632 ) , .A2( us12_n697 ) , .A1( us12_n724 ) );
  AOI21_X1 us12_U417 (.ZN( us12_n478 ) , .B2( us12_n697 ) , .A( us12_n749 ) , .B1( us12_n779 ) );
  NOR2_X1 us12_U418 (.A2( us12_n697 ) , .A1( us12_n780 ) , .ZN( us12_n820 ) );
  NOR2_X1 us12_U419 (.ZN( us12_n662 ) , .A2( us12_n697 ) , .A1( us12_n729 ) );
  AOI221_X1 us12_U42 (.A( us12_n781 ) , .ZN( us12_n798 ) , .C2( us12_n837 ) , .B2( us12_n838 ) , .B1( us12_n865 ) , .C1( us12_n866 ) );
  NOR2_X1 us12_U420 (.ZN( us12_n566 ) , .A2( us12_n697 ) , .A1( us12_n763 ) );
  NOR2_X1 us12_U421 (.ZN( us12_n600 ) , .A2( us12_n697 ) , .A1( us12_n784 ) );
  NOR2_X1 us12_U422 (.A2( us12_n697 ) , .ZN( us12_n716 ) , .A1( us12_n792 ) );
  NOR2_X1 us12_U423 (.ZN( us12_n594 ) , .A2( us12_n697 ) , .A1( us12_n728 ) );
  AOI21_X1 us12_U424 (.ZN( us12_n552 ) , .B1( us12_n669 ) , .A( us12_n697 ) , .B2( us12_n805 ) );
  NOR2_X1 us12_U425 (.ZN( us12_n541 ) , .A2( us12_n697 ) , .A1( us12_n699 ) );
  NOR2_X1 us12_U426 (.ZN( us12_n580 ) , .A2( us12_n697 ) , .A1( us12_n791 ) );
  NOR2_X1 us12_U427 (.A2( sa12_2 ) , .A1( sa12_3 ) , .ZN( us12_n472 ) );
  NOR2_X1 us12_U428 (.A2( sa12_3 ) , .ZN( us12_n455 ) , .A1( us12_n828 ) );
  INV_X1 us12_U429 (.A( sa12_3 ) , .ZN( us12_n829 ) );
  NOR4_X1 us12_U43 (.A4( us12_n793 ) , .A3( us12_n794 ) , .A2( us12_n795 ) , .A1( us12_n796 ) , .ZN( us12_n797 ) );
  OAI222_X1 us12_U430 (.ZN( us12_n505 ) , .C2( us12_n625 ) , .B2( us12_n647 ) , .B1( us12_n747 ) , .A2( us12_n748 ) , .C1( us12_n805 ) , .A1( us12_n806 ) );
  OAI222_X1 us12_U431 (.B2( us12_n747 ) , .B1( us12_n748 ) , .A2( us12_n749 ) , .ZN( us12_n757 ) , .C2( us12_n805 ) , .C1( us12_n814 ) , .A1( us12_n817 ) );
  NOR2_X1 us12_U432 (.ZN( us12_n748 ) , .A1( us12_n861 ) , .A2( us12_n862 ) );
  AND2_X1 us12_U433 (.ZN( us12_n438 ) , .A2( us12_n831 ) , .A1( us12_n854 ) );
  AND2_X1 us12_U434 (.ZN( us12_n439 ) , .A2( us12_n843 ) , .A1( us12_n861 ) );
  NOR3_X1 us12_U435 (.A1( us12_n438 ) , .A2( us12_n439 ) , .A3( us12_n576 ) , .ZN( us12_n587 ) );
  INV_X1 us12_U436 (.A( us12_n812 ) , .ZN( us12_n854 ) );
  NAND3_X1 us12_U437 (.ZN( sa11_sr_6 ) , .A3( us12_n797 ) , .A2( us12_n798 ) , .A1( us12_n799 ) );
  NAND3_X1 us12_U438 (.ZN( sa11_sr_5 ) , .A3( us12_n758 ) , .A2( us12_n759 ) , .A1( us12_n760 ) );
  NAND3_X1 us12_U439 (.ZN( sa11_sr_4 ) , .A3( us12_n738 ) , .A2( us12_n739 ) , .A1( us12_n740 ) );
  NOR4_X1 us12_U44 (.A4( us12_n776 ) , .A3( us12_n777 ) , .A1( us12_n778 ) , .ZN( us12_n799 ) , .A2( us12_n801 ) );
  NAND3_X1 us12_U440 (.A3( us12_n675 ) , .A2( us12_n676 ) , .A1( us12_n677 ) , .ZN( us12_n807 ) );
  NAND3_X1 us12_U441 (.ZN( us12_n638 ) , .A3( us12_n708 ) , .A2( us12_n724 ) , .A1( us12_n792 ) );
  NAND3_X1 us12_U442 (.A3( us12_n618 ) , .A2( us12_n619 ) , .A1( us12_n620 ) , .ZN( us12_n725 ) );
  NAND3_X1 us12_U443 (.A3( us12_n585 ) , .A2( us12_n586 ) , .A1( us12_n587 ) , .ZN( us12_n621 ) );
  NAND3_X1 us12_U444 (.ZN( us12_n565 ) , .A3( us12_n680 ) , .A2( us12_n750 ) , .A1( us12_n785 ) );
  NAND3_X1 us12_U445 (.A3( us12_n523 ) , .A2( us12_n524 ) , .A1( us12_n525 ) , .ZN( us12_n742 ) );
  NAND3_X1 us12_U446 (.A3( us12_n512 ) , .A1( us12_n513 ) , .ZN( us12_n608 ) , .A2( us12_n871 ) );
  NAND3_X1 us12_U447 (.A3( us12_n467 ) , .A2( us12_n468 ) , .A1( us12_n469 ) , .ZN( us12_n777 ) );
  INV_X1 us12_U448 (.A( us12_n803 ) , .ZN( us12_n843 ) );
  AOI21_X1 us12_U449 (.ZN( us12_n576 ) , .B2( us12_n724 ) , .B1( us12_n748 ) , .A( us12_n785 ) );
  NOR4_X1 us12_U45 (.A4( us12_n734 ) , .A3( us12_n735 ) , .A2( us12_n736 ) , .A1( us12_n737 ) , .ZN( us12_n738 ) );
  AOI211_X1 us12_U46 (.B( us12_n725 ) , .A( us12_n726 ) , .ZN( us12_n739 ) , .C1( us12_n843 ) , .C2( us12_n855 ) );
  NOR3_X1 us12_U47 (.A3( us12_n722 ) , .A1( us12_n723 ) , .ZN( us12_n740 ) , .A2( us12_n741 ) );
  NAND4_X1 us12_U48 (.ZN( sa11_sr_3 ) , .A4( us12_n704 ) , .A3( us12_n705 ) , .A2( us12_n706 ) , .A1( us12_n707 ) );
  NOR4_X1 us12_U49 (.A4( us12_n700 ) , .A3( us12_n701 ) , .A2( us12_n702 ) , .A1( us12_n703 ) , .ZN( us12_n704 ) );
  NAND2_X1 us12_U5 (.A2( us12_n448 ) , .A1( us12_n464 ) , .ZN( us12_n815 ) );
  AOI211_X1 us12_U50 (.B( us12_n694 ) , .A( us12_n695 ) , .ZN( us12_n705 ) , .C2( us12_n831 ) , .C1( us12_n851 ) );
  NOR2_X1 us12_U51 (.ZN( us12_n707 ) , .A2( us12_n776 ) , .A1( us12_n800 ) );
  NOR2_X1 us12_U52 (.ZN( us12_n804 ) , .A1( us12_n854 ) , .A2( us12_n861 ) );
  NAND4_X1 us12_U53 (.ZN( sa11_sr_0 ) , .A4( us12_n501 ) , .A3( us12_n502 ) , .A2( us12_n503 ) , .A1( us12_n504 ) );
  AOI221_X1 us12_U54 (.A( us12_n497 ) , .ZN( us12_n502 ) , .B2( us12_n843 ) , .C1( us12_n846 ) , .C2( us12_n860 ) , .B1( us12_n862 ) );
  NOR4_X1 us12_U55 (.A4( us12_n498 ) , .A3( us12_n499 ) , .A2( us12_n500 ) , .ZN( us12_n501 ) , .A1( us12_n527 ) );
  AOI211_X1 us12_U56 (.A( us12_n496 ) , .ZN( us12_n503 ) , .B( us12_n802 ) , .C2( us12_n839 ) , .C1( us12_n851 ) );
  NAND4_X1 us12_U57 (.ZN( sa11_sr_1 ) , .A4( us12_n595 ) , .A3( us12_n596 ) , .A2( us12_n597 ) , .A1( us12_n598 ) );
  AOI211_X1 us12_U58 (.B( us12_n589 ) , .A( us12_n590 ) , .ZN( us12_n596 ) , .C2( us12_n811 ) , .C1( us12_n833 ) );
  NOR4_X1 us12_U59 (.A4( us12_n591 ) , .A3( us12_n592 ) , .A2( us12_n593 ) , .A1( us12_n594 ) , .ZN( us12_n595 ) );
  NAND2_X1 us12_U6 (.A2( us12_n441 ) , .A1( us12_n452 ) , .ZN( us12_n791 ) );
  AOI211_X1 us12_U60 (.A( us12_n588 ) , .ZN( us12_n597 ) , .B( us12_n621 ) , .C1( us12_n845 ) , .C2( us12_n855 ) );
  NAND4_X1 us12_U61 (.ZN( sa11_sr_7 ) , .A4( us12_n822 ) , .A3( us12_n823 ) , .A2( us12_n824 ) , .A1( us12_n825 ) );
  NOR4_X1 us12_U62 (.A4( us12_n818 ) , .A3( us12_n819 ) , .A2( us12_n820 ) , .A1( us12_n821 ) , .ZN( us12_n822 ) );
  AOI222_X1 us12_U63 (.C2( us12_n809 ) , .B2( us12_n810 ) , .A2( us12_n811 ) , .ZN( us12_n823 ) , .C1( us12_n832 ) , .A1( us12_n839 ) , .B1( us12_n853 ) );
  AOI211_X1 us12_U64 (.B( us12_n807 ) , .A( us12_n808 ) , .ZN( us12_n824 ) , .C1( us12_n842 ) , .C2( us12_n850 ) );
  NAND4_X1 us12_U65 (.ZN( sa11_sr_2 ) , .A4( us12_n643 ) , .A3( us12_n644 ) , .A2( us12_n645 ) , .A1( us12_n646 ) );
  AOI222_X1 us12_U66 (.B2( us12_n638 ) , .ZN( us12_n644 ) , .B1( us12_n841 ) , .A1( us12_n842 ) , .C2( us12_n846 ) , .C1( us12_n863 ) , .A2( us12_n865 ) );
  NOR4_X1 us12_U67 (.A4( us12_n639 ) , .A3( us12_n640 ) , .A2( us12_n641 ) , .A1( us12_n642 ) , .ZN( us12_n643 ) );
  NOR3_X1 us12_U68 (.A2( us12_n607 ) , .A1( us12_n608 ) , .ZN( us12_n646 ) , .A3( us12_n722 ) );
  NAND4_X1 us12_U69 (.A4( us12_n603 ) , .A3( us12_n604 ) , .A2( us12_n605 ) , .A1( us12_n606 ) , .ZN( us12_n722 ) );
  NAND2_X1 us12_U7 (.A2( us12_n460 ) , .A1( us12_n465 ) , .ZN( us12_n780 ) );
  NOR3_X1 us12_U70 (.A1( us12_n599 ) , .ZN( us12_n604 ) , .A3( us12_n663 ) , .A2( us12_n770 ) );
  NOR4_X1 us12_U71 (.A3( us12_n600 ) , .A2( us12_n601 ) , .A1( us12_n602 ) , .ZN( us12_n603 ) , .A4( us12_n655 ) );
  AOI222_X1 us12_U72 (.ZN( us12_n606 ) , .A1( us12_n830 ) , .C2( us12_n837 ) , .B1( us12_n842 ) , .A2( us12_n856 ) , .B2( us12_n861 ) , .C1( us12_n868 ) );
  NOR4_X1 us12_U73 (.A4( us12_n514 ) , .A3( us12_n515 ) , .A2( us12_n516 ) , .A1( us12_n517 ) , .ZN( us12_n524 ) );
  AOI222_X1 us12_U74 (.ZN( us12_n525 ) , .A1( us12_n834 ) , .B2( us12_n837 ) , .C1( us12_n844 ) , .C2( us12_n850 ) , .A2( us12_n852 ) , .B1( us12_n866 ) );
  NOR4_X1 us12_U75 (.A3( us12_n521 ) , .A1( us12_n522 ) , .ZN( us12_n523 ) , .A2( us12_n673 ) , .A4( us12_n769 ) );
  NAND4_X1 us12_U76 (.A4( us12_n657 ) , .A3( us12_n658 ) , .A2( us12_n659 ) , .A1( us12_n660 ) , .ZN( us12_n800 ) );
  NOR3_X1 us12_U77 (.A3( us12_n648 ) , .A2( us12_n649 ) , .A1( us12_n650 ) , .ZN( us12_n659 ) );
  NOR3_X1 us12_U78 (.A3( us12_n651 ) , .A2( us12_n652 ) , .A1( us12_n653 ) , .ZN( us12_n658 ) );
  NOR3_X1 us12_U79 (.A3( us12_n654 ) , .A2( us12_n655 ) , .A1( us12_n656 ) , .ZN( us12_n657 ) );
  NOR3_X1 us12_U8 (.ZN( us12_n598 ) , .A1( us12_n608 ) , .A3( us12_n723 ) , .A2( us12_n742 ) );
  NAND4_X1 us12_U80 (.A4( us12_n560 ) , .A3( us12_n561 ) , .A2( us12_n562 ) , .A1( us12_n563 ) , .ZN( us12_n607 ) );
  NOR4_X1 us12_U81 (.A4( us12_n552 ) , .A3( us12_n553 ) , .A2( us12_n554 ) , .A1( us12_n555 ) , .ZN( us12_n562 ) );
  NOR4_X1 us12_U82 (.ZN( us12_n561 ) , .A1( us12_n653 ) , .A3( us12_n661 ) , .A4( us12_n685 ) , .A2( us12_n768 ) );
  NOR4_X1 us12_U83 (.A4( us12_n556 ) , .A3( us12_n557 ) , .A2( us12_n558 ) , .A1( us12_n559 ) , .ZN( us12_n560 ) );
  NAND4_X1 us12_U84 (.A4( us12_n772 ) , .A3( us12_n773 ) , .A2( us12_n774 ) , .A1( us12_n775 ) , .ZN( us12_n801 ) );
  NOR3_X1 us12_U85 (.A3( us12_n765 ) , .A2( us12_n766 ) , .A1( us12_n767 ) , .ZN( us12_n773 ) );
  NOR4_X1 us12_U86 (.A4( us12_n768 ) , .A3( us12_n769 ) , .A2( us12_n770 ) , .A1( us12_n771 ) , .ZN( us12_n772 ) );
  AOI222_X1 us12_U87 (.ZN( us12_n775 ) , .A1( us12_n830 ) , .C1( us12_n834 ) , .B2( us12_n841 ) , .A2( us12_n850 ) , .B1( us12_n861 ) , .C2( us12_n873 ) );
  NOR2_X1 us12_U88 (.ZN( us12_n625 ) , .A2( us12_n836 ) , .A1( us12_n839 ) );
  NOR2_X1 us12_U89 (.ZN( us12_n761 ) , .A1( us12_n833 ) , .A2( us12_n834 ) );
  NOR3_X1 us12_U9 (.A3( us12_n800 ) , .A2( us12_n801 ) , .A1( us12_n802 ) , .ZN( us12_n825 ) );
  AOI222_X1 us12_U90 (.ZN( us12_n513 ) , .C1( us12_n832 ) , .B2( us12_n837 ) , .A2( us12_n843 ) , .C2( us12_n862 ) , .B1( us12_n863 ) , .A1( us12_n866 ) );
  NOR4_X1 us12_U91 (.A4( us12_n509 ) , .A2( us12_n510 ) , .A1( us12_n511 ) , .ZN( us12_n512 ) , .A3( us12_n670 ) );
  INV_X1 us12_U92 (.A( us12_n505 ) , .ZN( us12_n871 ) );
  NAND4_X1 us12_U93 (.A4( us12_n456 ) , .A3( us12_n457 ) , .A2( us12_n458 ) , .A1( us12_n459 ) , .ZN( us12_n679 ) );
  NOR3_X1 us12_U94 (.ZN( us12_n457 ) , .A3( us12_n530 ) , .A1( us12_n555 ) , .A2( us12_n570 ) );
  AOI221_X1 us12_U95 (.A( us12_n450 ) , .ZN( us12_n459 ) , .C2( us12_n753 ) , .B1( us12_n832 ) , .C1( us12_n842 ) , .B2( us12_n861 ) );
  NOR4_X1 us12_U96 (.ZN( us12_n458 ) , .A2( us12_n509 ) , .A1( us12_n599 ) , .A4( us12_n628 ) , .A3( us12_n711 ) );
  NAND4_X1 us12_U97 (.A4( us12_n535 ) , .A3( us12_n536 ) , .A2( us12_n537 ) , .A1( us12_n538 ) , .ZN( us12_n622 ) );
  NOR4_X1 us12_U98 (.A4( us12_n526 ) , .A2( us12_n527 ) , .A1( us12_n528 ) , .ZN( us12_n538 ) , .A3( us12_n701 ) );
  NOR4_X1 us12_U99 (.A1( us12_n531 ) , .ZN( us12_n536 ) , .A2( us12_n654 ) , .A4( us12_n668 ) , .A3( us12_n765 ) );
  NOR3_X1 us31_U10 (.A3( us31_n621 ) , .A2( us31_n622 ) , .ZN( us31_n636 ) , .A1( us31_n725 ) );
  NOR4_X1 us31_U100 (.ZN( us31_n458 ) , .A2( us31_n509 ) , .A1( us31_n599 ) , .A4( us31_n628 ) , .A3( us31_n711 ) );
  NAND4_X1 us31_U101 (.A4( us31_n535 ) , .A3( us31_n536 ) , .A2( us31_n537 ) , .A1( us31_n538 ) , .ZN( us31_n622 ) );
  NOR4_X1 us31_U102 (.A4( us31_n526 ) , .A2( us31_n527 ) , .A1( us31_n528 ) , .ZN( us31_n538 ) , .A3( us31_n701 ) );
  NOR4_X1 us31_U103 (.A1( us31_n531 ) , .ZN( us31_n536 ) , .A2( us31_n654 ) , .A4( us31_n668 ) , .A3( us31_n765 ) );
  NOR4_X1 us31_U104 (.A4( us31_n529 ) , .A3( us31_n530 ) , .ZN( us31_n537 ) , .A2( us31_n684 ) , .A1( us31_n794 ) );
  NOR2_X1 us31_U105 (.ZN( us31_n647 ) , .A1( us31_n854 ) , .A2( us31_n868 ) );
  NAND4_X1 us31_U106 (.A4( us31_n548 ) , .A3( us31_n549 ) , .A2( us31_n550 ) , .A1( us31_n551 ) , .ZN( us31_n745 ) );
  NOR3_X1 us31_U107 (.ZN( us31_n549 ) , .A2( us31_n651 ) , .A1( us31_n667 ) , .A3( us31_n771 ) );
  AOI211_X1 us31_U108 (.B( us31_n539 ) , .A( us31_n540 ) , .ZN( us31_n551 ) , .C2( us31_n839 ) , .C1( us31_n851 ) );
  NOR4_X1 us31_U109 (.A4( us31_n541 ) , .A3( us31_n542 ) , .A2( us31_n543 ) , .ZN( us31_n550 ) , .A1( us31_n688 ) );
  NOR2_X1 us31_U11 (.A1( us31_n678 ) , .ZN( us31_n693 ) , .A2( us31_n807 ) );
  NAND4_X1 us31_U110 (.A4( us31_n479 ) , .A3( us31_n480 ) , .A2( us31_n481 ) , .A1( us31_n482 ) , .ZN( us31_n694 ) );
  NOR3_X1 us31_U111 (.ZN( us31_n480 ) , .A2( us31_n508 ) , .A3( us31_n601 ) , .A1( us31_n610 ) );
  AOI211_X1 us31_U112 (.B( us31_n477 ) , .A( us31_n478 ) , .ZN( us31_n482 ) , .C2( us31_n833 ) , .C1( us31_n861 ) );
  NOR4_X1 us31_U113 (.ZN( us31_n481 ) , .A3( us31_n532 ) , .A4( us31_n545 ) , .A2( us31_n567 ) , .A1( us31_n717 ) );
  NOR2_X1 us31_U114 (.ZN( us31_n686 ) , .A1( us31_n831 ) , .A2( us31_n832 ) );
  NAND4_X1 us31_U115 (.A4( us31_n485 ) , .A3( us31_n486 ) , .A2( us31_n487 ) , .A1( us31_n488 ) , .ZN( us31_n778 ) );
  NOR4_X1 us31_U116 (.A4( us31_n484 ) , .ZN( us31_n487 ) , .A1( us31_n566 ) , .A2( us31_n581 ) , .A3( us31_n602 ) );
  NOR4_X1 us31_U117 (.ZN( us31_n486 ) , .A1( us31_n507 ) , .A2( us31_n519 ) , .A4( us31_n546 ) , .A3( us31_n611 ) );
  NOR4_X1 us31_U118 (.ZN( us31_n485 ) , .A2( us31_n533 ) , .A1( us31_n558 ) , .A3( us31_n631 ) , .A4( us31_n718 ) );
  NAND4_X1 us31_U119 (.A4( us31_n691 ) , .A3( us31_n692 ) , .A1( us31_n693 ) , .ZN( us31_n776 ) , .A2( us31_n872 ) );
  NOR2_X1 us31_U12 (.ZN( us31_n495 ) , .A1( us31_n678 ) , .A2( us31_n694 ) );
  AOI221_X1 us31_U120 (.A( us31_n681 ) , .ZN( us31_n692 ) , .B2( us31_n840 ) , .C1( us31_n842 ) , .C2( us31_n862 ) , .B1( us31_n865 ) );
  INV_X1 us31_U121 (.A( us31_n679 ) , .ZN( us31_n872 ) );
  NOR4_X1 us31_U122 (.A4( us31_n687 ) , .A3( us31_n688 ) , .A2( us31_n689 ) , .A1( us31_n690 ) , .ZN( us31_n691 ) );
  NAND4_X1 us31_U123 (.A4( us31_n719 ) , .A3( us31_n720 ) , .A2( us31_n721 ) , .ZN( us31_n741 ) , .A1( us31_n857 ) );
  INV_X1 us31_U124 (.A( us31_n709 ) , .ZN( us31_n857 ) );
  AOI221_X1 us31_U125 (.A( us31_n710 ) , .ZN( us31_n721 ) , .C2( us31_n844 ) , .B2( us31_n845 ) , .C1( us31_n861 ) , .B1( us31_n862 ) );
  NOR4_X1 us31_U126 (.A4( us31_n715 ) , .A3( us31_n716 ) , .A2( us31_n717 ) , .A1( us31_n718 ) , .ZN( us31_n719 ) );
  NAND4_X1 us31_U127 (.A4( us31_n473 ) , .A3( us31_n474 ) , .A2( us31_n475 ) , .A1( us31_n476 ) , .ZN( us31_n678 ) );
  NOR4_X1 us31_U128 (.ZN( us31_n475 ) , .A1( us31_n531 ) , .A3( us31_n568 ) , .A4( us31_n600 ) , .A2( us31_n642 ) );
  NOR4_X1 us31_U129 (.ZN( us31_n473 ) , .A2( us31_n521 ) , .A4( us31_n594 ) , .A1( us31_n609 ) , .A3( us31_n629 ) );
  NOR3_X1 us31_U13 (.ZN( us31_n504 ) , .A2( us31_n679 ) , .A3( us31_n777 ) , .A1( us31_n876 ) );
  NOR4_X1 us31_U130 (.A4( us31_n470 ) , .ZN( us31_n476 ) , .A3( us31_n556 ) , .A1( us31_n735 ) , .A2( us31_n755 ) );
  NOR2_X1 us31_U131 (.ZN( us31_n733 ) , .A2( us31_n832 ) , .A1( us31_n845 ) );
  NOR2_X1 us31_U132 (.ZN( us31_n789 ) , .A2( us31_n862 ) , .A1( us31_n868 ) );
  NAND4_X1 us31_U133 (.A4( us31_n573 ) , .A3( us31_n574 ) , .A1( us31_n575 ) , .ZN( us31_n723 ) , .A2( us31_n874 ) );
  NOR4_X1 us31_U134 (.A4( us31_n569 ) , .A3( us31_n570 ) , .A2( us31_n571 ) , .A1( us31_n572 ) , .ZN( us31_n573 ) );
  AOI221_X1 us31_U135 (.A( us31_n564 ) , .C2( us31_n565 ) , .ZN( us31_n574 ) , .B2( us31_n845 ) , .B1( us31_n852 ) , .C1( us31_n853 ) );
  NOR2_X1 us31_U136 (.ZN( us31_n575 ) , .A1( us31_n622 ) , .A2( us31_n745 ) );
  NAND4_X1 us31_U137 (.A4( us31_n633 ) , .A3( us31_n634 ) , .A2( us31_n635 ) , .A1( us31_n636 ) , .ZN( us31_n743 ) );
  AOI211_X1 us31_U138 (.B( us31_n623 ) , .A( us31_n624 ) , .ZN( us31_n635 ) , .C2( us31_n836 ) , .C1( us31_n863 ) );
  NOR4_X1 us31_U139 (.A4( us31_n629 ) , .A3( us31_n630 ) , .A2( us31_n631 ) , .A1( us31_n632 ) , .ZN( us31_n633 ) );
  INV_X1 us31_U14 (.A( us31_n706 ) , .ZN( us31_n876 ) );
  NOR4_X1 us31_U140 (.A4( us31_n626 ) , .A3( us31_n627 ) , .A2( us31_n628 ) , .ZN( us31_n634 ) , .A1( us31_n664 ) );
  NAND4_X1 us31_U141 (.A4( us31_n493 ) , .A3( us31_n494 ) , .A1( us31_n495 ) , .ZN( us31_n802 ) , .A2( us31_n867 ) );
  AOI221_X1 us31_U142 (.A( us31_n489 ) , .ZN( us31_n494 ) , .B2( us31_n836 ) , .C2( us31_n841 ) , .C1( us31_n851 ) , .B1( us31_n860 ) );
  INV_X1 us31_U143 (.A( us31_n778 ) , .ZN( us31_n867 ) );
  NOR4_X1 us31_U144 (.A2( us31_n491 ) , .A1( us31_n492 ) , .ZN( us31_n493 ) , .A3( us31_n580 ) , .A4( us31_n612 ) );
  NOR4_X1 us31_U145 (.A4( us31_n734 ) , .A3( us31_n735 ) , .A2( us31_n736 ) , .A1( us31_n737 ) , .ZN( us31_n738 ) );
  AOI211_X1 us31_U146 (.B( us31_n725 ) , .A( us31_n726 ) , .ZN( us31_n739 ) , .C1( us31_n843 ) , .C2( us31_n855 ) );
  NOR3_X1 us31_U147 (.A3( us31_n722 ) , .A1( us31_n723 ) , .ZN( us31_n740 ) , .A2( us31_n741 ) );
  INV_X1 us31_U148 (.A( us31_n762 ) , .ZN( us31_n830 ) );
  INV_X1 us31_U149 (.A( us31_n697 ) , .ZN( us31_n838 ) );
  INV_X1 us31_U15 (.A( us31_n607 ) , .ZN( us31_n874 ) );
  OR4_X1 us31_U150 (.A4( us31_n566 ) , .A3( us31_n567 ) , .A2( us31_n568 ) , .ZN( us31_n572 ) , .A1( us31_n665 ) );
  OR4_X1 us31_U151 (.A4( us31_n682 ) , .A3( us31_n683 ) , .A2( us31_n684 ) , .A1( us31_n685 ) , .ZN( us31_n690 ) );
  OR4_X1 us31_U152 (.ZN( us31_n466 ) , .A4( us31_n518 ) , .A3( us31_n529 ) , .A2( us31_n578 ) , .A1( us31_n712 ) );
  OR4_X1 us31_U153 (.A4( us31_n518 ) , .A2( us31_n519 ) , .A1( us31_n520 ) , .ZN( us31_n522 ) , .A3( us31_n821 ) );
  OR4_X1 us31_U154 (.ZN( us31_n492 ) , .A4( us31_n534 ) , .A2( us31_n547 ) , .A1( us31_n559 ) , .A3( us31_n632 ) );
  OR4_X1 us31_U155 (.A4( us31_n580 ) , .A3( us31_n581 ) , .A2( us31_n582 ) , .A1( us31_n583 ) , .ZN( us31_n584 ) );
  NAND2_X1 us31_U156 (.ZN( us31_n613 ) , .A2( us31_n837 ) , .A1( us31_n873 ) );
  OR3_X1 us31_U157 (.A3( us31_n506 ) , .A2( us31_n507 ) , .A1( us31_n508 ) , .ZN( us31_n511 ) );
  INV_X1 us31_U158 (.A( us31_n463 ) , .ZN( us31_n864 ) );
  OAI21_X1 us31_U159 (.ZN( us31_n463 ) , .B1( us31_n809 ) , .A( us31_n834 ) , .B2( us31_n851 ) );
  INV_X1 us31_U16 (.A( us31_n680 ) , .ZN( us31_n840 ) );
  INV_X1 us31_U160 (.A( us31_n754 ) , .ZN( us31_n869 ) );
  OAI21_X1 us31_U161 (.B1( us31_n753 ) , .ZN( us31_n754 ) , .A( us31_n845 ) , .B2( us31_n868 ) );
  INV_X1 us31_U162 (.A( us31_n672 ) , .ZN( us31_n859 ) );
  AOI21_X1 us31_U163 (.A( us31_n670 ) , .B1( us31_n671 ) , .ZN( us31_n672 ) , .B2( us31_n856 ) );
  OAI222_X1 us31_U164 (.B2( us31_n747 ) , .B1( us31_n748 ) , .A2( us31_n749 ) , .ZN( us31_n757 ) , .C2( us31_n805 ) , .C1( us31_n814 ) , .A1( us31_n817 ) );
  OAI222_X1 us31_U165 (.ZN( us31_n505 ) , .C2( us31_n625 ) , .B2( us31_n647 ) , .B1( us31_n747 ) , .A2( us31_n748 ) , .C1( us31_n805 ) , .A1( us31_n806 ) );
  OAI222_X1 us31_U166 (.B2( us31_n708 ) , .ZN( us31_n709 ) , .C2( us31_n724 ) , .B1( us31_n747 ) , .A1( us31_n806 ) , .C1( us31_n814 ) , .A2( us31_n815 ) );
  NAND2_X1 us31_U167 (.A1( us31_n447 ) , .A2( us31_n465 ) , .ZN( us31_n749 ) );
  AOI22_X1 us31_U168 (.ZN( us31_n696 ) , .A1( us31_n830 ) , .B2( us31_n843 ) , .A2( us31_n865 ) , .B1( us31_n868 ) );
  AOI22_X1 us31_U169 (.A2( us31_n782 ) , .ZN( us31_n783 ) , .B2( us31_n831 ) , .A1( us31_n834 ) , .B1( us31_n863 ) );
  NOR4_X1 us31_U17 (.A4( us31_n445 ) , .A3( us31_n446 ) , .A2( us31_n516 ) , .A1( us31_n541 ) , .ZN( us31_n706 ) );
  INV_X1 us31_U170 (.A( us31_n730 ) , .ZN( us31_n839 ) );
  AOI221_X1 us31_U171 (.A( us31_n764 ) , .ZN( us31_n774 ) , .C2( us31_n810 ) , .B2( us31_n835 ) , .C1( us31_n855 ) , .B1( us31_n866 ) );
  AOI21_X1 us31_U172 (.B2( us31_n763 ) , .ZN( us31_n764 ) , .A( us31_n788 ) , .B1( us31_n792 ) );
  INV_X1 us31_U173 (.A( us31_n761 ) , .ZN( us31_n835 ) );
  AOI221_X1 us31_U174 (.A( us31_n483 ) , .ZN( us31_n488 ) , .B1( us31_n831 ) , .C2( us31_n844 ) , .C1( us31_n852 ) , .B2( us31_n862 ) );
  OAI22_X1 us31_U175 (.ZN( us31_n483 ) , .A1( us31_n708 ) , .B2( us31_n785 ) , .A2( us31_n806 ) , .B1( us31_n812 ) );
  INV_X1 us31_U176 (.A( us31_n790 ) , .ZN( us31_n832 ) );
  NAND2_X1 us31_U177 (.A1( us31_n451 ) , .A2( us31_n453 ) , .ZN( us31_n762 ) );
  AOI211_X1 us31_U178 (.A( us31_n637 ) , .ZN( us31_n645 ) , .B( us31_n743 ) , .C2( us31_n839 ) , .C1( us31_n854 ) );
  OAI22_X1 us31_U179 (.ZN( us31_n637 ) , .A1( us31_n699 ) , .B2( us31_n728 ) , .A2( us31_n762 ) , .B1( us31_n816 ) );
  OR3_X1 us31_U18 (.ZN( us31_n446 ) , .A1( us31_n528 ) , .A3( us31_n577 ) , .A2( us31_n875 ) );
  INV_X1 us31_U180 (.A( us31_n786 ) , .ZN( us31_n862 ) );
  OAI221_X1 us31_U181 (.A( us31_n727 ) , .C2( us31_n728 ) , .B2( us31_n729 ) , .B1( us31_n730 ) , .ZN( us31_n737 ) , .C1( us31_n817 ) );
  AOI22_X1 us31_U182 (.ZN( us31_n727 ) , .B1( us31_n832 ) , .A2( us31_n838 ) , .A1( us31_n863 ) , .B2( us31_n866 ) );
  OAI22_X1 us31_U183 (.ZN( us31_n710 ) , .A2( us31_n728 ) , .B2( us31_n729 ) , .A1( us31_n744 ) , .B1( us31_n813 ) );
  INV_X1 us31_U184 (.A( us31_n816 ) , .ZN( us31_n831 ) );
  OAI22_X1 us31_U185 (.ZN( us31_n624 ) , .B1( us31_n669 ) , .B2( us31_n747 ) , .A1( us31_n815 ) , .A2( us31_n816 ) );
  INV_X1 us31_U186 (.A( us31_n744 ) , .ZN( us31_n837 ) );
  INV_X1 us31_U187 (.A( us31_n788 ) , .ZN( us31_n845 ) );
  OAI22_X1 us31_U188 (.B2( us31_n779 ) , .B1( us31_n780 ) , .ZN( us31_n781 ) , .A2( us31_n814 ) , .A1( us31_n815 ) );
  OAI22_X1 us31_U189 (.A1( us31_n724 ) , .ZN( us31_n726 ) , .B2( us31_n750 ) , .B1( us31_n812 ) , .A2( us31_n816 ) );
  OR4_X1 us31_U19 (.A4( us31_n442 ) , .A2( us31_n443 ) , .A1( us31_n444 ) , .ZN( us31_n445 ) , .A3( us31_n553 ) );
  INV_X1 us31_U190 (.A( us31_n805 ) , .ZN( us31_n860 ) );
  INV_X1 us31_U191 (.A( us31_n814 ) , .ZN( us31_n833 ) );
  INV_X1 us31_U192 (.A( us31_n669 ) , .ZN( us31_n865 ) );
  OAI22_X1 us31_U193 (.B2( us31_n744 ) , .ZN( us31_n746 ) , .A2( us31_n762 ) , .B1( us31_n780 ) , .A1( us31_n792 ) );
  OAI22_X1 us31_U194 (.ZN( us31_n496 ) , .A2( us31_n744 ) , .A1( us31_n780 ) , .B1( us31_n791 ) , .B2( us31_n806 ) );
  OAI22_X1 us31_U195 (.B2( us31_n803 ) , .B1( us31_n804 ) , .A2( us31_n805 ) , .A1( us31_n806 ) , .ZN( us31_n808 ) );
  OAI22_X1 us31_U196 (.ZN( us31_n489 ) , .A1( us31_n724 ) , .B2( us31_n728 ) , .B1( us31_n730 ) , .A2( us31_n779 ) );
  OAI22_X1 us31_U197 (.ZN( us31_n695 ) , .A2( us31_n730 ) , .A1( us31_n780 ) , .B1( us31_n791 ) , .B2( us31_n817 ) );
  OAI22_X1 us31_U198 (.B1( us31_n490 ) , .ZN( us31_n491 ) , .A1( us31_n686 ) , .A2( us31_n763 ) , .B2( us31_n817 ) );
  NOR3_X1 us31_U199 (.ZN( us31_n490 ) , .A1( us31_n782 ) , .A2( us31_n850 ) , .A3( us31_n863 ) );
  INV_X1 us31_U20 (.A( us31_n613 ) , .ZN( us31_n875 ) );
  INV_X1 us31_U200 (.A( us31_n750 ) , .ZN( us31_n842 ) );
  NOR2_X1 us31_U201 (.ZN( us31_n715 ) , .A1( us31_n805 ) , .A2( us31_n817 ) );
  NOR2_X1 us31_U202 (.A2( us31_n744 ) , .ZN( us31_n755 ) , .A1( us31_n805 ) );
  NOR2_X1 us31_U203 (.ZN( us31_n735 ) , .A2( us31_n803 ) , .A1( us31_n805 ) );
  NOR2_X1 us31_U204 (.ZN( us31_n546 ) , .A2( us31_n780 ) , .A1( us31_n814 ) );
  NOR2_X1 us31_U205 (.ZN( us31_n577 ) , .A2( us31_n699 ) , .A1( us31_n814 ) );
  NOR2_X1 us31_U206 (.ZN( us31_n718 ) , .A2( us31_n724 ) , .A1( us31_n744 ) );
  NOR2_X1 us31_U207 (.ZN( us31_n532 ) , .A2( us31_n749 ) , .A1( us31_n750 ) );
  NOR2_X1 us31_U208 (.ZN( us31_n615 ) , .A1( us31_n785 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U209 (.ZN( us31_n629 ) , .A2( us31_n728 ) , .A1( us31_n785 ) );
  INV_X1 us31_U21 (.A( us31_n749 ) , .ZN( us31_n863 ) );
  NOR2_X1 us31_U210 (.ZN( us31_n611 ) , .A2( us31_n780 ) , .A1( us31_n806 ) );
  NOR2_X1 us31_U211 (.ZN( us31_n652 ) , .A1( us31_n669 ) , .A2( us31_n814 ) );
  NOR2_X1 us31_U212 (.A1( us31_n669 ) , .ZN( us31_n673 ) , .A2( us31_n744 ) );
  NOR2_X1 us31_U213 (.ZN( us31_n602 ) , .A1( us31_n669 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U214 (.A1( us31_n669 ) , .ZN( us31_n688 ) , .A2( us31_n816 ) );
  NOR2_X1 us31_U215 (.ZN( us31_n628 ) , .A2( us31_n669 ) , .A1( us31_n785 ) );
  INV_X1 us31_U216 (.A( us31_n747 ) , .ZN( us31_n834 ) );
  NOR2_X1 us31_U217 (.A1( us31_n669 ) , .ZN( us31_n766 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U218 (.A2( us31_n744 ) , .ZN( us31_n769 ) , .A1( us31_n812 ) );
  NOR2_X1 us31_U219 (.ZN( us31_n527 ) , .A1( us31_n669 ) , .A2( us31_n779 ) );
  AOI222_X1 us31_U22 (.ZN( us31_n605 ) , .B2( us31_n671 ) , .B1( us31_n753 ) , .C2( us31_n831 ) , .A1( us31_n833 ) , .A2( us31_n862 ) , .C1( us31_n863 ) );
  NOR2_X1 us31_U220 (.ZN( us31_n531 ) , .A2( us31_n780 ) , .A1( us31_n816 ) );
  INV_X1 us31_U221 (.A( us31_n792 ) , .ZN( us31_n851 ) );
  NOR2_X1 us31_U222 (.A2( us31_n708 ) , .A1( us31_n750 ) , .ZN( us31_n771 ) );
  NOR2_X1 us31_U223 (.ZN( us31_n599 ) , .A2( us31_n791 ) , .A1( us31_n816 ) );
  NOR2_X1 us31_U224 (.ZN( us31_n601 ) , .A2( us31_n780 ) , .A1( us31_n803 ) );
  NOR2_X1 us31_U225 (.A1( us31_n699 ) , .ZN( us31_n768 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U226 (.ZN( us31_n541 ) , .A2( us31_n697 ) , .A1( us31_n699 ) );
  NOR2_X1 us31_U227 (.ZN( us31_n667 ) , .A1( us31_n750 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U228 (.ZN( us31_n555 ) , .A1( us31_n750 ) , .A2( us31_n791 ) );
  NOR2_X1 us31_U229 (.ZN( us31_n508 ) , .A2( us31_n780 ) , .A1( us31_n785 ) );
  AOI222_X1 us31_U23 (.ZN( us31_n563 ) , .B1( us31_n830 ) , .C1( us31_n841 ) , .A2( us31_n843 ) , .A1( us31_n854 ) , .B2( us31_n863 ) , .C2( us31_n873 ) );
  NOR2_X1 us31_U230 (.ZN( us31_n543 ) , .A2( us31_n708 ) , .A1( us31_n785 ) );
  NOR2_X1 us31_U231 (.ZN( us31_n528 ) , .A2( us31_n724 ) , .A1( us31_n803 ) );
  NOR2_X1 us31_U232 (.ZN( us31_n664 ) , .A1( us31_n785 ) , .A2( us31_n791 ) );
  NOR2_X1 us31_U233 (.ZN( us31_n556 ) , .A1( us31_n762 ) , .A2( us31_n805 ) );
  INV_X1 us31_U234 (.A( us31_n806 ) , .ZN( us31_n841 ) );
  OAI22_X1 us31_U235 (.B1( us31_n440 ) , .ZN( us31_n444 ) , .A2( us31_n728 ) , .A1( us31_n744 ) , .B2( us31_n749 ) );
  NOR3_X1 us31_U236 (.ZN( us31_n440 ) , .A2( us31_n836 ) , .A3( us31_n837 ) , .A1( us31_n846 ) );
  NOR2_X1 us31_U237 (.ZN( us31_n507 ) , .A1( us31_n812 ) , .A2( us31_n817 ) );
  NOR2_X1 us31_U238 (.ZN( us31_n557 ) , .A1( us31_n792 ) , .A2( us31_n814 ) );
  NOR2_X1 us31_U239 (.ZN( us31_n545 ) , .A1( us31_n749 ) , .A2( us31_n814 ) );
  AOI222_X1 us31_U24 (.ZN( us31_n660 ) , .A2( us31_n839 ) , .B1( us31_n841 ) , .C2( us31_n845 ) , .A1( us31_n860 ) , .C1( us31_n863 ) , .B2( us31_n870 ) );
  OAI22_X1 us31_U240 (.B2( us31_n750 ) , .B1( us31_n751 ) , .A1( us31_n752 ) , .ZN( us31_n756 ) , .A2( us31_n806 ) );
  NOR2_X1 us31_U241 (.ZN( us31_n751 ) , .A2( us31_n852 ) , .A1( us31_n860 ) );
  NOR3_X1 us31_U242 (.ZN( us31_n752 ) , .A2( us31_n853 ) , .A1( us31_n863 ) , .A3( us31_n865 ) );
  NOR2_X1 us31_U243 (.ZN( us31_n544 ) , .A2( us31_n785 ) , .A1( us31_n792 ) );
  NOR2_X1 us31_U244 (.ZN( us31_n530 ) , .A2( us31_n744 ) , .A1( us31_n792 ) );
  NOR2_X1 us31_U245 (.ZN( us31_n509 ) , .A1( us31_n729 ) , .A2( us31_n779 ) );
  NOR2_X1 us31_U246 (.ZN( us31_n570 ) , .A1( us31_n728 ) , .A2( us31_n806 ) );
  NOR2_X1 us31_U247 (.ZN( us31_n666 ) , .A1( us31_n728 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U248 (.ZN( us31_n631 ) , .A1( us31_n724 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U249 (.ZN( us31_n614 ) , .A1( us31_n762 ) , .A2( us31_n812 ) );
  INV_X1 us31_U25 (.A( us31_n647 ) , .ZN( us31_n870 ) );
  NOR2_X1 us31_U250 (.A1( us31_n749 ) , .ZN( us31_n767 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U251 (.ZN( us31_n654 ) , .A1( us31_n728 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U252 (.ZN( us31_n516 ) , .A1( us31_n708 ) , .A2( us31_n744 ) );
  NOR2_X1 us31_U253 (.ZN( us31_n670 ) , .A1( us31_n790 ) , .A2( us31_n805 ) );
  NOR2_X1 us31_U254 (.ZN( us31_n558 ) , .A1( us31_n708 ) , .A2( us31_n816 ) );
  INV_X1 us31_U255 (.A( us31_n763 ) , .ZN( us31_n866 ) );
  NOR2_X1 us31_U256 (.ZN( us31_n663 ) , .A1( us31_n729 ) , .A2( us31_n785 ) );
  NOR2_X1 us31_U257 (.A2( us31_n697 ) , .ZN( us31_n716 ) , .A1( us31_n792 ) );
  NOR2_X1 us31_U258 (.ZN( us31_n517 ) , .A1( us31_n708 ) , .A2( us31_n803 ) );
  NOR2_X1 us31_U259 (.ZN( us31_n521 ) , .A1( us31_n790 ) , .A2( us31_n812 ) );
  NOR4_X1 us31_U26 (.A4( us31_n544 ) , .A3( us31_n545 ) , .A2( us31_n546 ) , .A1( us31_n547 ) , .ZN( us31_n548 ) );
  NOR2_X1 us31_U260 (.ZN( us31_n630 ) , .A1( us31_n747 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U261 (.ZN( us31_n655 ) , .A1( us31_n790 ) , .A2( us31_n815 ) );
  AOI21_X1 us31_U262 (.ZN( us31_n552 ) , .B1( us31_n669 ) , .A( us31_n697 ) , .B2( us31_n805 ) );
  NOR2_X1 us31_U263 (.ZN( us31_n668 ) , .A2( us31_n708 ) , .A1( us31_n790 ) );
  NOR2_X1 us31_U264 (.ZN( us31_n594 ) , .A2( us31_n697 ) , .A1( us31_n728 ) );
  NOR2_X1 us31_U265 (.ZN( us31_n542 ) , .A1( us31_n762 ) , .A2( us31_n791 ) );
  NOR2_X1 us31_U266 (.ZN( us31_n656 ) , .A1( us31_n747 ) , .A2( us31_n780 ) );
  NOR2_X1 us31_U267 (.ZN( us31_n609 ) , .A2( us31_n724 ) , .A1( us31_n817 ) );
  AOI21_X1 us31_U268 (.B1( us31_n625 ) , .ZN( us31_n627 ) , .A( us31_n763 ) , .B2( us31_n814 ) );
  NOR2_X1 us31_U269 (.ZN( us31_n661 ) , .A1( us31_n729 ) , .A2( us31_n790 ) );
  NOR4_X1 us31_U27 (.ZN( us31_n479 ) , .A1( us31_n520 ) , .A4( us31_n557 ) , .A3( us31_n582 ) , .A2( us31_n630 ) );
  NOR2_X1 us31_U270 (.ZN( us31_n642 ) , .A2( us31_n788 ) , .A1( us31_n791 ) );
  AOI21_X1 us31_U271 (.ZN( us31_n650 ) , .A( us31_n779 ) , .B1( us31_n792 ) , .B2( us31_n805 ) );
  AOI21_X1 us31_U272 (.ZN( us31_n626 ) , .B2( us31_n669 ) , .A( us31_n790 ) , .B1( us31_n791 ) );
  AOI21_X1 us31_U273 (.A( us31_n815 ) , .B2( us31_n816 ) , .B1( us31_n817 ) , .ZN( us31_n818 ) );
  NOR2_X1 us31_U274 (.ZN( us31_n579 ) , .A2( us31_n708 ) , .A1( us31_n730 ) );
  NOR2_X1 us31_U275 (.ZN( us31_n533 ) , .A2( us31_n724 ) , .A1( us31_n730 ) );
  AOI21_X1 us31_U276 (.A( us31_n812 ) , .B2( us31_n813 ) , .B1( us31_n814 ) , .ZN( us31_n819 ) );
  NOR2_X1 us31_U277 (.A2( us31_n708 ) , .A1( us31_n762 ) , .ZN( us31_n794 ) );
  NOR2_X1 us31_U278 (.A2( us31_n697 ) , .A1( us31_n780 ) , .ZN( us31_n820 ) );
  AOI21_X1 us31_U279 (.ZN( us31_n499 ) , .B1( us31_n680 ) , .A( us31_n812 ) , .B2( us31_n816 ) );
  NOR4_X1 us31_U28 (.ZN( us31_n456 ) , .A2( us31_n517 ) , .A1( us31_n543 ) , .A3( us31_n579 ) , .A4( us31_n615 ) );
  NOR2_X1 us31_U280 (.ZN( us31_n520 ) , .A2( us31_n708 ) , .A1( us31_n814 ) );
  AOI21_X1 us31_U281 (.ZN( us31_n477 ) , .A( us31_n669 ) , .B1( us31_n750 ) , .B2( us31_n806 ) );
  NOR2_X1 us31_U282 (.ZN( us31_n582 ) , .A1( us31_n744 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U283 (.ZN( us31_n662 ) , .A2( us31_n697 ) , .A1( us31_n729 ) );
  AOI21_X1 us31_U284 (.ZN( us31_n593 ) , .B1( us31_n750 ) , .A( us31_n792 ) , .B2( us31_n813 ) );
  AOI21_X1 us31_U285 (.ZN( us31_n515 ) , .A( us31_n729 ) , .B1( us31_n750 ) , .B2( us31_n803 ) );
  AOI21_X1 us31_U286 (.ZN( us31_n510 ) , .B2( us31_n669 ) , .A( us31_n730 ) , .B1( us31_n815 ) );
  NOR2_X1 us31_U287 (.ZN( us31_n506 ) , .A2( us31_n728 ) , .A1( us31_n762 ) );
  NOR2_X1 us31_U288 (.A1( us31_n697 ) , .ZN( us31_n770 ) , .A2( us31_n815 ) );
  NOR2_X1 us31_U289 (.ZN( us31_n519 ) , .A2( us31_n699 ) , .A1( us31_n816 ) );
  NOR4_X1 us31_U29 (.A4( us31_n532 ) , .A3( us31_n533 ) , .A2( us31_n534 ) , .ZN( us31_n535 ) , .A1( us31_n820 ) );
  NOR2_X1 us31_U290 (.ZN( us31_n581 ) , .A1( us31_n669 ) , .A2( us31_n788 ) );
  NOR2_X1 us31_U291 (.ZN( us31_n559 ) , .A2( us31_n791 ) , .A1( us31_n803 ) );
  AOI21_X1 us31_U292 (.B1( us31_n699 ) , .ZN( us31_n700 ) , .A( us31_n732 ) , .B2( us31_n763 ) );
  AOI21_X1 us31_U293 (.ZN( us31_n591 ) , .B2( us31_n763 ) , .A( us31_n785 ) , .B1( us31_n812 ) );
  INV_X1 us31_U294 (.A( us31_n813 ) , .ZN( us31_n836 ) );
  NOR2_X1 us31_U295 (.ZN( us31_n683 ) , .A2( us31_n699 ) , .A1( us31_n803 ) );
  AOI21_X1 us31_U296 (.ZN( us31_n589 ) , .B2( us31_n699 ) , .B1( us31_n815 ) , .A( us31_n817 ) );
  AOI21_X1 us31_U297 (.ZN( us31_n539 ) , .B2( us31_n812 ) , .A( us31_n814 ) , .B1( us31_n815 ) );
  INV_X1 us31_U298 (.A( us31_n728 ) , .ZN( us31_n852 ) );
  AOI21_X1 us31_U299 (.ZN( us31_n540 ) , .A( us31_n763 ) , .B2( us31_n779 ) , .B1( us31_n817 ) );
  NAND2_X1 us31_U3 (.A1( us31_n449 ) , .A2( us31_n460 ) , .ZN( us31_n792 ) );
  NOR4_X1 us31_U30 (.ZN( us31_n474 ) , .A1( us31_n506 ) , .A3( us31_n544 ) , .A2( us31_n583 ) , .A4( us31_n716 ) );
  INV_X1 us31_U300 (.A( us31_n791 ) , .ZN( us31_n873 ) );
  AOI21_X1 us31_U301 (.ZN( us31_n498 ) , .A( us31_n724 ) , .B2( us31_n762 ) , .B1( us31_n814 ) );
  AOI21_X1 us31_U302 (.ZN( us31_n649 ) , .B1( us31_n729 ) , .B2( us31_n763 ) , .A( us31_n813 ) );
  NOR2_X1 us31_U303 (.ZN( us31_n547 ) , .A1( us31_n699 ) , .A2( us31_n744 ) );
  NOR2_X1 us31_U304 (.ZN( us31_n566 ) , .A2( us31_n697 ) , .A1( us31_n763 ) );
  AOI21_X1 us31_U305 (.ZN( us31_n569 ) , .B1( us31_n750 ) , .B2( us31_n762 ) , .A( us31_n780 ) );
  AOI21_X1 us31_U306 (.ZN( us31_n571 ) , .B2( us31_n697 ) , .B1( us31_n806 ) , .A( us31_n812 ) );
  AOI21_X1 us31_U307 (.ZN( us31_n640 ) , .B2( us31_n747 ) , .A( us31_n792 ) , .B1( us31_n803 ) );
  INV_X1 us31_U308 (.A( us31_n699 ) , .ZN( us31_n853 ) );
  AOI21_X1 us31_U309 (.ZN( us31_n514 ) , .A( us31_n779 ) , .B2( us31_n792 ) , .B1( us31_n812 ) );
  AOI221_X1 us31_U31 (.A( us31_n713 ) , .B2( us31_n714 ) , .ZN( us31_n720 ) , .C1( us31_n832 ) , .B1( us31_n839 ) , .C2( us31_n863 ) );
  AOI21_X1 us31_U310 (.ZN( us31_n639 ) , .B2( us31_n749 ) , .A( us31_n788 ) , .B1( us31_n812 ) );
  NAND2_X1 us31_U311 (.ZN( us31_n753 ) , .A1( us31_n763 ) , .A2( us31_n805 ) );
  NOR2_X1 us31_U312 (.ZN( us31_n665 ) , .A1( us31_n780 ) , .A2( us31_n813 ) );
  INV_X1 us31_U313 (.A( us31_n729 ) , .ZN( us31_n868 ) );
  NOR2_X1 us31_U314 (.ZN( us31_n685 ) , .A1( us31_n729 ) , .A2( us31_n816 ) );
  AOI21_X1 us31_U315 (.ZN( us31_n564 ) , .B1( us31_n724 ) , .A( us31_n779 ) , .B2( us31_n791 ) );
  AOI21_X1 us31_U316 (.ZN( us31_n497 ) , .A( us31_n779 ) , .B2( us31_n791 ) , .B1( us31_n804 ) );
  AOI21_X1 us31_U317 (.ZN( us31_n689 ) , .B2( us31_n749 ) , .B1( us31_n763 ) , .A( us31_n806 ) );
  AOI21_X1 us31_U318 (.ZN( us31_n450 ) , .B2( us31_n792 ) , .A( us31_n803 ) , .B1( us31_n815 ) );
  NOR2_X1 us31_U319 (.ZN( us31_n567 ) , .A1( us31_n747 ) , .A2( us31_n805 ) );
  OR2_X1 us31_U32 (.A2( us31_n711 ) , .A1( us31_n712 ) , .ZN( us31_n713 ) );
  NOR2_X1 us31_U320 (.ZN( us31_n529 ) , .A1( us31_n708 ) , .A2( us31_n779 ) );
  NOR2_X1 us31_U321 (.ZN( us31_n578 ) , .A1( us31_n708 ) , .A2( us31_n813 ) );
  AOI21_X1 us31_U322 (.ZN( us31_n478 ) , .B2( us31_n697 ) , .A( us31_n749 ) , .B1( us31_n779 ) );
  AOI21_X1 us31_U323 (.A( us31_n790 ) , .B2( us31_n791 ) , .B1( us31_n792 ) , .ZN( us31_n793 ) );
  NOR2_X1 us31_U324 (.ZN( us31_n684 ) , .A1( us31_n791 ) , .A2( us31_n813 ) );
  AOI21_X1 us31_U325 (.A( us31_n733 ) , .ZN( us31_n734 ) , .B2( us31_n780 ) , .B1( us31_n792 ) );
  NOR2_X1 us31_U326 (.A2( us31_n813 ) , .A1( us31_n815 ) , .ZN( us31_n821 ) );
  NOR2_X1 us31_U327 (.ZN( us31_n711 ) , .A1( us31_n762 ) , .A2( us31_n763 ) );
  AOI21_X1 us31_U328 (.ZN( us31_n641 ) , .B1( us31_n680 ) , .A( us31_n791 ) , .B2( us31_n817 ) );
  NOR2_X1 us31_U329 (.ZN( us31_n580 ) , .A2( us31_n697 ) , .A1( us31_n791 ) );
  NOR2_X1 us31_U33 (.ZN( us31_n680 ) , .A2( us31_n834 ) , .A1( us31_n839 ) );
  NOR2_X1 us31_U330 (.ZN( us31_n583 ) , .A1( us31_n792 ) , .A2( us31_n817 ) );
  NOR2_X1 us31_U331 (.ZN( us31_n534 ) , .A1( us31_n724 ) , .A2( us31_n788 ) );
  NOR2_X1 us31_U332 (.ZN( us31_n632 ) , .A2( us31_n697 ) , .A1( us31_n724 ) );
  NOR2_X1 us31_U333 (.ZN( us31_n682 ) , .A2( us31_n708 ) , .A1( us31_n817 ) );
  AOI21_X1 us31_U334 (.B1( us31_n686 ) , .ZN( us31_n687 ) , .A( us31_n728 ) , .B2( us31_n761 ) );
  INV_X1 us31_U335 (.A( us31_n815 ) , .ZN( us31_n855 ) );
  AOI21_X1 us31_U336 (.ZN( us31_n442 ) , .A( us31_n699 ) , .B1( us31_n733 ) , .B2( us31_n750 ) );
  NOR2_X1 us31_U337 (.ZN( us31_n568 ) , .A1( us31_n729 ) , .A2( us31_n762 ) );
  INV_X1 us31_U338 (.A( us31_n780 ) , .ZN( us31_n850 ) );
  INV_X1 us31_U339 (.A( us31_n785 ) , .ZN( us31_n846 ) );
  AOI222_X1 us31_U34 (.ZN( us31_n469 ) , .B1( us31_n832 ) , .A1( us31_n839 ) , .C1( us31_n842 ) , .C2( us31_n851 ) , .A2( us31_n855 ) , .B2( us31_n865 ) );
  NAND2_X1 us31_U340 (.A2( us31_n762 ) , .A1( us31_n806 ) , .ZN( us31_n810 ) );
  AOI21_X1 us31_U341 (.ZN( us31_n443 ) , .B1( us31_n789 ) , .B2( us31_n791 ) , .A( us31_n814 ) );
  NAND2_X1 us31_U342 (.ZN( us31_n671 ) , .A1( us31_n806 ) , .A2( us31_n816 ) );
  NOR2_X1 us31_U343 (.ZN( us31_n484 ) , .A1( us31_n788 ) , .A2( us31_n805 ) );
  NOR2_X1 us31_U344 (.ZN( us31_n470 ) , .A2( us31_n779 ) , .A1( us31_n815 ) );
  NOR2_X1 us31_U345 (.ZN( us31_n712 ) , .A2( us31_n724 ) , .A1( us31_n790 ) );
  OAI21_X1 us31_U346 (.A( us31_n787 ) , .B2( us31_n788 ) , .B1( us31_n789 ) , .ZN( us31_n795 ) );
  OAI21_X1 us31_U347 (.ZN( us31_n787 ) , .A( us31_n839 ) , .B1( us31_n863 ) , .B2( us31_n873 ) );
  NOR2_X1 us31_U348 (.ZN( us31_n526 ) , .A1( us31_n724 ) , .A2( us31_n750 ) );
  NAND2_X1 us31_U349 (.A1( us31_n699 ) , .A2( us31_n729 ) , .ZN( us31_n782 ) );
  NOR4_X1 us31_U35 (.A1( us31_n466 ) , .ZN( us31_n467 ) , .A4( us31_n542 ) , .A2( us31_n554 ) , .A3( us31_n614 ) );
  NOR2_X1 us31_U350 (.ZN( us31_n518 ) , .A1( us31_n708 ) , .A2( us31_n788 ) );
  OAI21_X1 us31_U351 (.A( us31_n698 ) , .ZN( us31_n702 ) , .B2( us31_n750 ) , .B1( us31_n804 ) );
  OAI21_X1 us31_U352 (.ZN( us31_n698 ) , .B2( us31_n833 ) , .B1( us31_n838 ) , .A( us31_n860 ) );
  INV_X1 us31_U353 (.A( us31_n817 ) , .ZN( us31_n844 ) );
  OAI21_X1 us31_U354 (.A( us31_n731 ) , .B1( us31_n732 ) , .ZN( us31_n736 ) , .B2( us31_n805 ) );
  OAI21_X1 us31_U355 (.ZN( us31_n731 ) , .A( us31_n833 ) , .B2( us31_n852 ) , .B1( us31_n873 ) );
  NAND2_X1 us31_U356 (.ZN( us31_n714 ) , .A1( us31_n728 ) , .A2( us31_n780 ) );
  INV_X1 us31_U357 (.A( us31_n724 ) , .ZN( us31_n856 ) );
  AND2_X1 us31_U358 (.ZN( us31_n732 ) , .A1( us31_n779 ) , .A2( us31_n785 ) );
  NAND2_X1 us31_U359 (.A1( us31_n447 ) , .A2( us31_n449 ) , .ZN( us31_n805 ) );
  AOI221_X1 us31_U36 (.ZN( us31_n468 ) , .C2( us31_n714 ) , .B2( us31_n831 ) , .C1( us31_n845 ) , .B1( us31_n860 ) , .A( us31_n864 ) );
  NAND2_X1 us31_U360 (.A1( us31_n451 ) , .A2( us31_n454 ) , .ZN( us31_n814 ) );
  NAND2_X1 us31_U361 (.A1( us31_n452 ) , .A2( us31_n465 ) , .ZN( us31_n669 ) );
  NAND2_X1 us31_U362 (.A1( us31_n455 ) , .A2( us31_n462 ) , .ZN( us31_n750 ) );
  NAND2_X1 us31_U363 (.A2( us31_n453 ) , .A1( us31_n455 ) , .ZN( us31_n806 ) );
  NAND2_X1 us31_U364 (.A1( us31_n451 ) , .A2( us31_n471 ) , .ZN( us31_n816 ) );
  NAND2_X1 us31_U365 (.A1( us31_n454 ) , .A2( us31_n461 ) , .ZN( us31_n813 ) );
  NAND2_X1 us31_U366 (.A1( us31_n455 ) , .A2( us31_n471 ) , .ZN( us31_n803 ) );
  NAND2_X1 us31_U367 (.A1( us31_n453 ) , .A2( us31_n461 ) , .ZN( us31_n744 ) );
  NAND2_X1 us31_U368 (.A1( us31_n453 ) , .A2( us31_n472 ) , .ZN( us31_n785 ) );
  NAND2_X1 us31_U369 (.A2( us31_n454 ) , .A1( us31_n472 ) , .ZN( us31_n779 ) );
  NOR4_X1 us31_U37 (.A4( us31_n577 ) , .A3( us31_n578 ) , .A2( us31_n579 ) , .ZN( us31_n586 ) , .A1( us31_n683 ) );
  NAND2_X1 us31_U370 (.A2( us31_n464 ) , .A1( us31_n465 ) , .ZN( us31_n812 ) );
  NAND2_X1 us31_U371 (.A1( us31_n441 ) , .A2( us31_n460 ) , .ZN( us31_n699 ) );
  NAND2_X1 us31_U372 (.A2( us31_n449 ) , .A1( us31_n452 ) , .ZN( us31_n763 ) );
  NAND2_X1 us31_U373 (.A2( us31_n461 ) , .A1( us31_n462 ) , .ZN( us31_n747 ) );
  NAND2_X1 us31_U374 (.A1( us31_n462 ) , .A2( us31_n472 ) , .ZN( us31_n788 ) );
  NOR2_X1 us31_U375 (.ZN( us31_n465 ) , .A2( us31_n847 ) , .A1( us31_n848 ) );
  NOR2_X1 us31_U376 (.ZN( us31_n453 ) , .A1( us31_n826 ) , .A2( us31_n827 ) );
  NOR2_X1 us31_U377 (.ZN( us31_n451 ) , .A1( us31_n828 ) , .A2( us31_n829 ) );
  NAND2_X1 us31_U378 (.A1( us31_n451 ) , .A2( us31_n462 ) , .ZN( us31_n790 ) );
  NAND2_X1 us31_U379 (.A2( us31_n441 ) , .A1( us31_n447 ) , .ZN( us31_n784 ) );
  NOR4_X1 us31_U38 (.A1( us31_n584 ) , .ZN( us31_n585 ) , .A3( us31_n652 ) , .A2( us31_n662 ) , .A4( us31_n767 ) );
  NAND2_X1 us31_U380 (.A2( us31_n454 ) , .A1( us31_n455 ) , .ZN( us31_n730 ) );
  NAND2_X2 us31_U381 (.A1( us31_n449 ) , .A2( us31_n464 ) , .ZN( us31_n724 ) );
  NAND2_X2 us31_U382 (.A2( us31_n460 ) , .A1( us31_n465 ) , .ZN( us31_n780 ) );
  NOR2_X1 us31_U383 (.ZN( us31_n447 ) , .A2( us31_n849 ) , .A1( us31_n858 ) );
  NAND2_X1 us31_U384 (.A1( us31_n447 ) , .A2( us31_n448 ) , .ZN( us31_n786 ) );
  NAND2_X1 us31_U385 (.A2( us31_n448 ) , .A1( us31_n460 ) , .ZN( us31_n728 ) );
  NAND2_X1 us31_U386 (.A2( us31_n448 ) , .A1( us31_n452 ) , .ZN( us31_n729 ) );
  NOR2_X1 us31_U387 (.A2( sa31_5 ) , .ZN( us31_n448 ) , .A1( us31_n847 ) );
  NOR2_X1 us31_U388 (.A2( sa31_7 ) , .ZN( us31_n460 ) , .A1( us31_n849 ) );
  NOR2_X1 us31_U389 (.A2( sa31_6 ) , .A1( sa31_7 ) , .ZN( us31_n464 ) );
  NOR4_X1 us31_U39 (.ZN( us31_n620 ) , .A1( us31_n656 ) , .A3( us31_n666 ) , .A4( us31_n682 ) , .A2( us31_n766 ) );
  NOR2_X1 us31_U390 (.A2( sa31_4 ) , .ZN( us31_n449 ) , .A1( us31_n848 ) );
  NOR2_X1 us31_U391 (.A2( sa31_4 ) , .A1( sa31_5 ) , .ZN( us31_n441 ) );
  NOR2_X1 us31_U392 (.A2( sa31_6 ) , .ZN( us31_n452 ) , .A1( us31_n858 ) );
  NOR2_X1 us31_U393 (.A2( sa31_2 ) , .A1( sa31_3 ) , .ZN( us31_n472 ) );
  NOR2_X1 us31_U394 (.A2( sa31_1 ) , .ZN( us31_n471 ) , .A1( us31_n826 ) );
  NOR2_X1 us31_U395 (.A2( sa31_0 ) , .ZN( us31_n454 ) , .A1( us31_n827 ) );
  NOR2_X1 us31_U396 (.A2( sa31_0 ) , .A1( sa31_1 ) , .ZN( us31_n462 ) );
  NOR2_X1 us31_U397 (.A2( sa31_3 ) , .ZN( us31_n455 ) , .A1( us31_n828 ) );
  NOR2_X1 us31_U398 (.A2( sa31_2 ) , .ZN( us31_n461 ) , .A1( us31_n829 ) );
  INV_X1 us31_U399 (.A( sa31_4 ) , .ZN( us31_n847 ) );
  NAND2_X1 us31_U4 (.A2( us31_n448 ) , .A1( us31_n464 ) , .ZN( us31_n815 ) );
  NOR4_X1 us31_U40 (.A4( us31_n609 ) , .A3( us31_n610 ) , .A2( us31_n611 ) , .A1( us31_n612 ) , .ZN( us31_n619 ) );
  INV_X1 us31_U400 (.A( sa31_6 ) , .ZN( us31_n849 ) );
  INV_X1 us31_U401 (.A( sa31_3 ) , .ZN( us31_n829 ) );
  INV_X1 us31_U402 (.A( sa31_1 ) , .ZN( us31_n827 ) );
  INV_X1 us31_U403 (.A( sa31_0 ) , .ZN( us31_n826 ) );
  INV_X1 us31_U404 (.A( sa31_2 ) , .ZN( us31_n828 ) );
  INV_X1 us31_U405 (.A( sa31_5 ) , .ZN( us31_n848 ) );
  INV_X1 us31_U406 (.A( sa31_7 ) , .ZN( us31_n858 ) );
  NAND2_X1 us31_U407 (.A2( us31_n461 ) , .A1( us31_n471 ) , .ZN( us31_n697 ) );
  OAI22_X1 us31_U408 (.ZN( us31_n588 ) , .A2( us31_n747 ) , .B2( us31_n762 ) , .A1( us31_n763 ) , .B1( us31_n784 ) );
  AOI21_X1 us31_U409 (.ZN( us31_n592 ) , .B1( us31_n728 ) , .B2( us31_n784 ) , .A( us31_n790 ) );
  NOR4_X1 us31_U41 (.A4( us31_n614 ) , .A3( us31_n615 ) , .A2( us31_n616 ) , .A1( us31_n617 ) , .ZN( us31_n618 ) );
  NAND2_X1 us31_U410 (.A1( us31_n729 ) , .A2( us31_n784 ) , .ZN( us31_n811 ) );
  AOI21_X1 us31_U411 (.ZN( us31_n623 ) , .B1( us31_n699 ) , .A( us31_n779 ) , .B2( us31_n784 ) );
  OAI22_X1 us31_U412 (.ZN( us31_n681 ) , .A1( us31_n699 ) , .A2( us31_n730 ) , .B2( us31_n784 ) , .B1( us31_n817 ) );
  AOI21_X1 us31_U413 (.ZN( us31_n648 ) , .A( us31_n762 ) , .B2( us31_n784 ) , .B1( us31_n792 ) );
  OAI21_X1 us31_U414 (.A( us31_n613 ) , .ZN( us31_n616 ) , .B1( us31_n625 ) , .B2( us31_n784 ) );
  OAI222_X1 us31_U415 (.A2( us31_n669 ) , .ZN( us31_n674 ) , .B1( us31_n747 ) , .B2( us31_n784 ) , .C2( us31_n788 ) , .C1( us31_n815 ) , .A1( us31_n817 ) );
  NOR2_X1 us31_U416 (.ZN( us31_n610 ) , .A1( us31_n784 ) , .A2( us31_n816 ) );
  NOR2_X1 us31_U417 (.ZN( us31_n651 ) , .A1( us31_n784 ) , .A2( us31_n788 ) );
  NOR2_X1 us31_U418 (.ZN( us31_n553 ) , .A2( us31_n744 ) , .A1( us31_n784 ) );
  NOR2_X1 us31_U419 (.ZN( us31_n600 ) , .A2( us31_n697 ) , .A1( us31_n784 ) );
  NOR4_X1 us31_U42 (.A4( us31_n514 ) , .A3( us31_n515 ) , .A2( us31_n516 ) , .A1( us31_n517 ) , .ZN( us31_n524 ) );
  INV_X1 us31_U420 (.A( us31_n784 ) , .ZN( us31_n861 ) );
  AND2_X1 us31_U421 (.ZN( us31_n438 ) , .A2( us31_n831 ) , .A1( us31_n854 ) );
  AND2_X1 us31_U422 (.ZN( us31_n439 ) , .A2( us31_n843 ) , .A1( us31_n861 ) );
  NOR3_X1 us31_U423 (.A1( us31_n438 ) , .A2( us31_n439 ) , .A3( us31_n576 ) , .ZN( us31_n587 ) );
  INV_X1 us31_U424 (.A( us31_n812 ) , .ZN( us31_n854 ) );
  INV_X1 us31_U425 (.A( us31_n803 ) , .ZN( us31_n843 ) );
  AOI21_X1 us31_U426 (.ZN( us31_n576 ) , .B2( us31_n724 ) , .B1( us31_n748 ) , .A( us31_n785 ) );
  OAI221_X1 us31_U427 (.A( us31_n783 ) , .C2( us31_n784 ) , .B2( us31_n785 ) , .B1( us31_n786 ) , .ZN( us31_n796 ) , .C1( us31_n813 ) );
  AOI21_X1 us31_U428 (.ZN( us31_n500 ) , .A( us31_n697 ) , .B1( us31_n708 ) , .B2( us31_n786 ) );
  OAI221_X1 us31_U429 (.A( us31_n696 ) , .ZN( us31_n703 ) , .C2( us31_n784 ) , .C1( us31_n785 ) , .B1( us31_n786 ) , .B2( us31_n806 ) );
  AOI222_X1 us31_U43 (.ZN( us31_n525 ) , .A1( us31_n834 ) , .B2( us31_n837 ) , .C1( us31_n844 ) , .C2( us31_n850 ) , .A2( us31_n852 ) , .B1( us31_n866 ) );
  OAI22_X1 us31_U430 (.ZN( us31_n590 ) , .B1( us31_n730 ) , .B2( us31_n749 ) , .A2( us31_n786 ) , .A1( us31_n803 ) );
  NAND2_X1 us31_U431 (.A2( us31_n749 ) , .A1( us31_n786 ) , .ZN( us31_n809 ) );
  NOR2_X1 us31_U432 (.ZN( us31_n612 ) , .A1( us31_n779 ) , .A2( us31_n786 ) );
  OAI222_X1 us31_U433 (.ZN( us31_n617 ) , .B1( us31_n697 ) , .C1( us31_n724 ) , .C2( us31_n747 ) , .B2( us31_n786 ) , .A2( us31_n792 ) , .A1( us31_n816 ) );
  NOR2_X1 us31_U434 (.ZN( us31_n653 ) , .A1( us31_n762 ) , .A2( us31_n786 ) );
  NOR2_X1 us31_U435 (.ZN( us31_n554 ) , .A1( us31_n786 ) , .A2( us31_n813 ) );
  NOR2_X1 us31_U436 (.ZN( us31_n717 ) , .A2( us31_n744 ) , .A1( us31_n786 ) );
  NAND3_X1 us31_U437 (.ZN( sa32_sr_6 ) , .A3( us31_n797 ) , .A2( us31_n798 ) , .A1( us31_n799 ) );
  NAND3_X1 us31_U438 (.ZN( sa32_sr_5 ) , .A3( us31_n758 ) , .A2( us31_n759 ) , .A1( us31_n760 ) );
  NAND3_X1 us31_U439 (.ZN( sa32_sr_4 ) , .A3( us31_n738 ) , .A2( us31_n739 ) , .A1( us31_n740 ) );
  NOR4_X1 us31_U44 (.A3( us31_n521 ) , .A1( us31_n522 ) , .ZN( us31_n523 ) , .A2( us31_n673 ) , .A4( us31_n769 ) );
  NAND3_X1 us31_U440 (.A3( us31_n675 ) , .A2( us31_n676 ) , .A1( us31_n677 ) , .ZN( us31_n807 ) );
  NAND3_X1 us31_U441 (.ZN( us31_n638 ) , .A3( us31_n708 ) , .A2( us31_n724 ) , .A1( us31_n792 ) );
  NAND3_X1 us31_U442 (.A3( us31_n618 ) , .A2( us31_n619 ) , .A1( us31_n620 ) , .ZN( us31_n725 ) );
  NAND3_X1 us31_U443 (.A3( us31_n585 ) , .A2( us31_n586 ) , .A1( us31_n587 ) , .ZN( us31_n621 ) );
  NAND3_X1 us31_U444 (.ZN( us31_n565 ) , .A3( us31_n680 ) , .A2( us31_n750 ) , .A1( us31_n785 ) );
  NAND3_X1 us31_U445 (.A3( us31_n523 ) , .A2( us31_n524 ) , .A1( us31_n525 ) , .ZN( us31_n742 ) );
  NAND3_X1 us31_U446 (.A3( us31_n512 ) , .A1( us31_n513 ) , .ZN( us31_n608 ) , .A2( us31_n871 ) );
  NAND3_X1 us31_U447 (.A3( us31_n467 ) , .A2( us31_n468 ) , .A1( us31_n469 ) , .ZN( us31_n777 ) );
  NOR2_X1 us31_U448 (.ZN( us31_n701 ) , .A2( us31_n786 ) , .A1( us31_n817 ) );
  NOR2_X1 us31_U449 (.A1( us31_n730 ) , .ZN( us31_n765 ) , .A2( us31_n786 ) );
  AOI221_X1 us31_U45 (.A( us31_n781 ) , .ZN( us31_n798 ) , .C2( us31_n837 ) , .B2( us31_n838 ) , .B1( us31_n865 ) , .C1( us31_n866 ) );
  NOR4_X1 us31_U46 (.A4( us31_n793 ) , .A3( us31_n794 ) , .A2( us31_n795 ) , .A1( us31_n796 ) , .ZN( us31_n797 ) );
  NOR4_X1 us31_U47 (.A4( us31_n776 ) , .A3( us31_n777 ) , .A1( us31_n778 ) , .ZN( us31_n799 ) , .A2( us31_n801 ) );
  NOR4_X1 us31_U48 (.A3( us31_n755 ) , .A2( us31_n756 ) , .A1( us31_n757 ) , .ZN( us31_n758 ) , .A4( us31_n869 ) );
  AOI211_X1 us31_U49 (.B( us31_n745 ) , .A( us31_n746 ) , .ZN( us31_n759 ) , .C1( us31_n832 ) , .C2( us31_n853 ) );
  NAND2_X1 us31_U5 (.A1( us31_n441 ) , .A2( us31_n464 ) , .ZN( us31_n708 ) );
  NOR3_X1 us31_U50 (.A3( us31_n741 ) , .A2( us31_n742 ) , .A1( us31_n743 ) , .ZN( us31_n760 ) );
  NAND4_X1 us31_U51 (.ZN( sa32_sr_3 ) , .A4( us31_n704 ) , .A3( us31_n705 ) , .A2( us31_n706 ) , .A1( us31_n707 ) );
  NOR4_X1 us31_U52 (.A4( us31_n700 ) , .A3( us31_n701 ) , .A2( us31_n702 ) , .A1( us31_n703 ) , .ZN( us31_n704 ) );
  AOI211_X1 us31_U53 (.B( us31_n694 ) , .A( us31_n695 ) , .ZN( us31_n705 ) , .C2( us31_n831 ) , .C1( us31_n851 ) );
  NOR2_X1 us31_U54 (.ZN( us31_n707 ) , .A2( us31_n776 ) , .A1( us31_n800 ) );
  NOR2_X1 us31_U55 (.ZN( us31_n804 ) , .A1( us31_n854 ) , .A2( us31_n861 ) );
  NAND4_X1 us31_U56 (.ZN( sa32_sr_7 ) , .A4( us31_n822 ) , .A3( us31_n823 ) , .A2( us31_n824 ) , .A1( us31_n825 ) );
  NOR4_X1 us31_U57 (.A4( us31_n818 ) , .A3( us31_n819 ) , .A2( us31_n820 ) , .A1( us31_n821 ) , .ZN( us31_n822 ) );
  AOI222_X1 us31_U58 (.C2( us31_n809 ) , .B2( us31_n810 ) , .A2( us31_n811 ) , .ZN( us31_n823 ) , .C1( us31_n832 ) , .A1( us31_n839 ) , .B1( us31_n853 ) );
  AOI211_X1 us31_U59 (.B( us31_n807 ) , .A( us31_n808 ) , .ZN( us31_n824 ) , .C1( us31_n842 ) , .C2( us31_n850 ) );
  NAND2_X1 us31_U6 (.A2( us31_n441 ) , .A1( us31_n452 ) , .ZN( us31_n791 ) );
  NAND4_X1 us31_U60 (.ZN( sa32_sr_0 ) , .A4( us31_n501 ) , .A3( us31_n502 ) , .A2( us31_n503 ) , .A1( us31_n504 ) );
  AOI221_X1 us31_U61 (.A( us31_n497 ) , .ZN( us31_n502 ) , .B2( us31_n843 ) , .C1( us31_n846 ) , .C2( us31_n860 ) , .B1( us31_n862 ) );
  NOR4_X1 us31_U62 (.A4( us31_n498 ) , .A3( us31_n499 ) , .A2( us31_n500 ) , .ZN( us31_n501 ) , .A1( us31_n527 ) );
  AOI211_X1 us31_U63 (.A( us31_n496 ) , .ZN( us31_n503 ) , .B( us31_n802 ) , .C2( us31_n839 ) , .C1( us31_n851 ) );
  NAND4_X1 us31_U64 (.ZN( sa32_sr_1 ) , .A4( us31_n595 ) , .A3( us31_n596 ) , .A2( us31_n597 ) , .A1( us31_n598 ) );
  NOR4_X1 us31_U65 (.A4( us31_n591 ) , .A3( us31_n592 ) , .A2( us31_n593 ) , .A1( us31_n594 ) , .ZN( us31_n595 ) );
  AOI211_X1 us31_U66 (.B( us31_n589 ) , .A( us31_n590 ) , .ZN( us31_n596 ) , .C2( us31_n811 ) , .C1( us31_n833 ) );
  AOI211_X1 us31_U67 (.A( us31_n588 ) , .ZN( us31_n597 ) , .B( us31_n621 ) , .C1( us31_n845 ) , .C2( us31_n855 ) );
  NAND4_X1 us31_U68 (.ZN( sa32_sr_2 ) , .A4( us31_n643 ) , .A3( us31_n644 ) , .A2( us31_n645 ) , .A1( us31_n646 ) );
  AOI222_X1 us31_U69 (.B2( us31_n638 ) , .ZN( us31_n644 ) , .B1( us31_n841 ) , .A1( us31_n842 ) , .C2( us31_n846 ) , .C1( us31_n863 ) , .A2( us31_n865 ) );
  NAND2_X1 us31_U7 (.A2( us31_n471 ) , .A1( us31_n472 ) , .ZN( us31_n817 ) );
  NOR4_X1 us31_U70 (.A4( us31_n639 ) , .A3( us31_n640 ) , .A2( us31_n641 ) , .A1( us31_n642 ) , .ZN( us31_n643 ) );
  NOR3_X1 us31_U71 (.A2( us31_n607 ) , .A1( us31_n608 ) , .ZN( us31_n646 ) , .A3( us31_n722 ) );
  NOR2_X1 us31_U72 (.ZN( us31_n748 ) , .A1( us31_n861 ) , .A2( us31_n862 ) );
  NOR2_X1 us31_U73 (.ZN( us31_n625 ) , .A2( us31_n836 ) , .A1( us31_n839 ) );
  NAND4_X1 us31_U74 (.A4( us31_n603 ) , .A3( us31_n604 ) , .A2( us31_n605 ) , .A1( us31_n606 ) , .ZN( us31_n722 ) );
  NOR3_X1 us31_U75 (.A1( us31_n599 ) , .ZN( us31_n604 ) , .A3( us31_n663 ) , .A2( us31_n770 ) );
  NOR4_X1 us31_U76 (.A3( us31_n600 ) , .A2( us31_n601 ) , .A1( us31_n602 ) , .ZN( us31_n603 ) , .A4( us31_n655 ) );
  AOI222_X1 us31_U77 (.ZN( us31_n606 ) , .A1( us31_n830 ) , .C2( us31_n837 ) , .B1( us31_n842 ) , .A2( us31_n856 ) , .B2( us31_n861 ) , .C1( us31_n868 ) );
  NAND4_X1 us31_U78 (.A4( us31_n657 ) , .A3( us31_n658 ) , .A2( us31_n659 ) , .A1( us31_n660 ) , .ZN( us31_n800 ) );
  NOR3_X1 us31_U79 (.A3( us31_n648 ) , .A2( us31_n649 ) , .A1( us31_n650 ) , .ZN( us31_n659 ) );
  NOR3_X1 us31_U8 (.ZN( us31_n598 ) , .A1( us31_n608 ) , .A3( us31_n723 ) , .A2( us31_n742 ) );
  NOR3_X1 us31_U80 (.A3( us31_n651 ) , .A2( us31_n652 ) , .A1( us31_n653 ) , .ZN( us31_n658 ) );
  NOR3_X1 us31_U81 (.A3( us31_n654 ) , .A2( us31_n655 ) , .A1( us31_n656 ) , .ZN( us31_n657 ) );
  NAND4_X1 us31_U82 (.A4( us31_n560 ) , .A3( us31_n561 ) , .A2( us31_n562 ) , .A1( us31_n563 ) , .ZN( us31_n607 ) );
  NOR4_X1 us31_U83 (.ZN( us31_n561 ) , .A1( us31_n653 ) , .A3( us31_n661 ) , .A4( us31_n685 ) , .A2( us31_n768 ) );
  NOR4_X1 us31_U84 (.A4( us31_n552 ) , .A3( us31_n553 ) , .A2( us31_n554 ) , .A1( us31_n555 ) , .ZN( us31_n562 ) );
  NOR4_X1 us31_U85 (.A4( us31_n556 ) , .A3( us31_n557 ) , .A2( us31_n558 ) , .A1( us31_n559 ) , .ZN( us31_n560 ) );
  NAND4_X1 us31_U86 (.A4( us31_n772 ) , .A3( us31_n773 ) , .A2( us31_n774 ) , .A1( us31_n775 ) , .ZN( us31_n801 ) );
  NOR3_X1 us31_U87 (.A3( us31_n765 ) , .A2( us31_n766 ) , .A1( us31_n767 ) , .ZN( us31_n773 ) );
  NOR4_X1 us31_U88 (.A4( us31_n768 ) , .A3( us31_n769 ) , .A2( us31_n770 ) , .A1( us31_n771 ) , .ZN( us31_n772 ) );
  AOI222_X1 us31_U89 (.ZN( us31_n775 ) , .A1( us31_n830 ) , .C1( us31_n834 ) , .B2( us31_n841 ) , .A2( us31_n850 ) , .B1( us31_n861 ) , .C2( us31_n873 ) );
  NOR3_X1 us31_U9 (.A3( us31_n800 ) , .A2( us31_n801 ) , .A1( us31_n802 ) , .ZN( us31_n825 ) );
  NOR4_X1 us31_U90 (.A4( us31_n661 ) , .A3( us31_n662 ) , .A2( us31_n663 ) , .A1( us31_n664 ) , .ZN( us31_n677 ) );
  NOR4_X1 us31_U91 (.A4( us31_n665 ) , .A3( us31_n666 ) , .A2( us31_n667 ) , .A1( us31_n668 ) , .ZN( us31_n676 ) );
  NOR4_X1 us31_U92 (.A3( us31_n673 ) , .A1( us31_n674 ) , .ZN( us31_n675 ) , .A4( us31_n715 ) , .A2( us31_n859 ) );
  NOR2_X1 us31_U93 (.ZN( us31_n761 ) , .A1( us31_n833 ) , .A2( us31_n834 ) );
  AOI222_X1 us31_U94 (.ZN( us31_n513 ) , .C1( us31_n832 ) , .B2( us31_n837 ) , .A2( us31_n843 ) , .C2( us31_n862 ) , .B1( us31_n863 ) , .A1( us31_n866 ) );
  NOR4_X1 us31_U95 (.A4( us31_n509 ) , .A2( us31_n510 ) , .A1( us31_n511 ) , .ZN( us31_n512 ) , .A3( us31_n670 ) );
  INV_X1 us31_U96 (.A( us31_n505 ) , .ZN( us31_n871 ) );
  NAND4_X1 us31_U97 (.A4( us31_n456 ) , .A3( us31_n457 ) , .A2( us31_n458 ) , .A1( us31_n459 ) , .ZN( us31_n679 ) );
  NOR3_X1 us31_U98 (.ZN( us31_n457 ) , .A3( us31_n530 ) , .A1( us31_n555 ) , .A2( us31_n570 ) );
  AOI221_X1 us31_U99 (.A( us31_n450 ) , .ZN( us31_n459 ) , .C2( us31_n753 ) , .B1( us31_n832 ) , .C1( us31_n842 ) , .B2( us31_n861 ) );
endmodule

