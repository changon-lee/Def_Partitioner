module des_des_die_6 ( u0_K12_34, u0_K12_35, u0_K12_36, u0_K12_39, u0_K12_40, u0_K12_48, u0_K13_45, u0_K13_46, u0_K13_48, 
       u0_L10_11, u0_L10_12, u0_L10_14, u0_L10_15, u0_L10_19, u0_L10_21, u0_L10_22, u0_L10_25, u0_L10_27, 
       u0_L10_29, u0_L10_3, u0_L10_32, u0_L10_4, u0_L10_5, u0_L10_7, u0_L10_8, u0_L11_15, u0_L11_17, 
       u0_L11_21, u0_L11_23, u0_L11_27, u0_L11_31, u0_L11_5, u0_L11_9, u0_L9_14, u0_L9_25, u0_L9_3, 
       u0_L9_8, u0_R10_1, u0_R10_16, u0_R10_17, u0_R10_18, u0_R10_19, u0_R10_20, u0_R10_21, u0_R10_22, 
       u0_R10_23, u0_R10_24, u0_R10_25, u0_R10_26, u0_R10_27, u0_R10_28, u0_R10_29, u0_R10_30, u0_R10_31, 
       u0_R10_32, u0_R11_1, u0_R11_2, u0_R11_28, u0_R11_29, u0_R11_3, u0_R11_30, u0_R11_31, u0_R11_32, 
       u0_R11_4, u0_R11_5, u0_R9_16, u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_20, u0_R9_21, u0_uk_K_r10_14, 
       u0_uk_K_r10_23, u0_uk_K_r10_28, u0_uk_K_r10_37, u0_uk_K_r10_42, u0_uk_K_r10_43, u0_uk_K_r10_44, u0_uk_K_r10_9, u0_uk_K_r11_19, u0_uk_K_r11_24, 
       u0_uk_K_r11_25, u0_uk_K_r11_26, u0_uk_K_r11_29, u0_uk_K_r11_4, u0_uk_K_r11_46, u0_uk_K_r11_48, u0_uk_K_r11_53, u0_uk_K_r9_0, u0_uk_K_r9_1, 
       u0_uk_K_r9_35, u0_uk_K_r9_9, u0_uk_n10, u0_uk_n100, u0_uk_n102, u0_uk_n106, u0_uk_n107, u0_uk_n109, u0_uk_n11, 
       u0_uk_n110, u0_uk_n117, u0_uk_n118, u0_uk_n119, u0_uk_n121, u0_uk_n126, u0_uk_n129, u0_uk_n131, u0_uk_n134, 
       u0_uk_n139, u0_uk_n140, u0_uk_n141, u0_uk_n142, u0_uk_n144, u0_uk_n145, u0_uk_n148, u0_uk_n151, u0_uk_n152, 
       u0_uk_n153, u0_uk_n154, u0_uk_n159, u0_uk_n161, u0_uk_n163, u0_uk_n167, u0_uk_n168, u0_uk_n171, u0_uk_n173, 
       u0_uk_n174, u0_uk_n178, u0_uk_n179, u0_uk_n180, u0_uk_n182, u0_uk_n184, u0_uk_n191, u0_uk_n192, u0_uk_n193, 
       u0_uk_n198, u0_uk_n203, u0_uk_n204, u0_uk_n207, u0_uk_n208, u0_uk_n211, u0_uk_n213, u0_uk_n214, u0_uk_n216, 
       u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n224, u0_uk_n238, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, 
       u0_uk_n31, u0_uk_n60, u0_uk_n83, u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n96, u0_uk_n99, u2_K10_32, 
       u2_K10_34, u2_K10_36, u2_K10_42, u2_K12_2, u2_K12_8, u2_K1_19, u2_K1_21, u2_K1_24, u2_K1_28, 
       u2_K1_37, u2_K1_40, u2_K1_43, u2_K1_45, u2_K1_46, u2_K2_34, u2_K2_35, u2_K2_36, u2_K2_40, 
       u2_K5_1, u2_K5_10, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_16, u2_K5_17, u2_K5_18, u2_K5_19, 
       u2_K5_21, u2_K5_23, u2_K5_24, u2_K5_25, u2_K5_26, u2_K5_28, u2_K5_3, u2_K5_5, u2_K5_6, 
       u2_K5_8, u2_K5_9, u2_K8_18, u2_K8_5, u2_K9_23, u2_K9_25, u2_K9_28, u2_K9_29, u2_L0_11, 
       u2_L0_12, u2_L0_19, u2_L0_22, u2_L0_29, u2_L0_32, u2_L0_4, u2_L0_7, u2_L10_13, u2_L10_17, 
       u2_L10_18, u2_L10_2, u2_L10_23, u2_L10_28, u2_L10_31, u2_L10_9, u2_L12_15, u2_L12_21, u2_L12_27, 
       u2_L12_5, u2_L3_1, u2_L3_10, u2_L3_13, u2_L3_14, u2_L3_16, u2_L3_17, u2_L3_18, u2_L3_2, 
       u2_L3_20, u2_L3_23, u2_L3_24, u2_L3_25, u2_L3_26, u2_L3_28, u2_L3_3, u2_L3_30, u2_L3_31, 
       u2_L3_6, u2_L3_8, u2_L3_9, u2_L6_16, u2_L6_17, u2_L6_23, u2_L6_24, u2_L6_30, u2_L6_31, 
       u2_L6_6, u2_L6_9, u2_L7_1, u2_L7_10, u2_L7_14, u2_L7_20, u2_L7_25, u2_L7_26, u2_L7_3, 
       u2_L7_8, u2_L8_11, u2_L8_12, u2_L8_19, u2_L8_22, u2_L8_29, u2_L8_32, u2_L8_4, u2_L8_7, 
       u2_R0_20, u2_R0_21, u2_R0_22, u2_R0_23, u2_R0_24, u2_R0_25, u2_R0_26, u2_R0_27, u2_R0_28, 
       u2_R0_29, u2_R10_1, u2_R10_2, u2_R10_3, u2_R10_32, u2_R10_4, u2_R10_5, u2_R10_6, u2_R10_7, 
       u2_R10_8, u2_R10_9, u2_R12_1, u2_R12_28, u2_R12_29, u2_R12_30, u2_R12_31, u2_R12_32, u2_R3_1, 
       u2_R3_10, u2_R3_11, u2_R3_12, u2_R3_13, u2_R3_14, u2_R3_15, u2_R3_16, u2_R3_17, u2_R3_18, 
       u2_R3_19, u2_R3_2, u2_R3_20, u2_R3_21, u2_R3_3, u2_R3_32, u2_R3_4, u2_R3_5, u2_R3_6, 
       u2_R3_7, u2_R3_8, u2_R3_9, u2_R6_1, u2_R6_10, u2_R6_11, u2_R6_12, u2_R6_13, u2_R6_2, 
       u2_R6_3, u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_8, u2_R6_9, u2_R7_12, u2_R7_13, u2_R7_14, 
       u2_R7_15, u2_R7_16, u2_R7_17, u2_R7_18, u2_R7_19, u2_R7_20, u2_R7_21, u2_R8_20, u2_R8_21, 
       u2_R8_22, u2_R8_23, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, u2_desIn_r_0, 
       u2_desIn_r_1, u2_desIn_r_11, u2_desIn_r_12, u2_desIn_r_16, u2_desIn_r_17, u2_desIn_r_18, u2_desIn_r_19, u2_desIn_r_20, u2_desIn_r_22, 
       u2_desIn_r_25, u2_desIn_r_26, u2_desIn_r_27, u2_desIn_r_28, u2_desIn_r_29, u2_desIn_r_3, u2_desIn_r_30, u2_desIn_r_32, u2_desIn_r_33, 
       u2_desIn_r_34, u2_desIn_r_35, u2_desIn_r_37, u2_desIn_r_38, u2_desIn_r_41, u2_desIn_r_42, u2_desIn_r_43, u2_desIn_r_44, u2_desIn_r_45, 
       u2_desIn_r_49, u2_desIn_r_51, u2_desIn_r_52, u2_desIn_r_53, u2_desIn_r_54, u2_desIn_r_56, u2_desIn_r_57, u2_desIn_r_59, u2_desIn_r_6, 
       u2_desIn_r_61, u2_desIn_r_62, u2_desIn_r_7, u2_desIn_r_8, u2_desIn_r_9, u2_key_r_0, u2_key_r_14, u2_key_r_16, u2_key_r_2, 
       u2_key_r_21, u2_key_r_22, u2_key_r_23, u2_key_r_25, u2_key_r_28, u2_key_r_29, u2_key_r_30, u2_key_r_31, u2_key_r_32, 
       u2_key_r_33, u2_key_r_35, u2_key_r_36, u2_key_r_37, u2_key_r_40, u2_key_r_42, u2_key_r_43, u2_key_r_44, u2_key_r_47, 
       u2_key_r_48, u2_key_r_51, u2_key_r_52, u2_key_r_55, u2_key_r_7, u2_key_r_9, u2_uk_K_r0_15, u2_uk_K_r0_31, u2_uk_K_r0_36, 
       u2_uk_K_r10_10, u2_uk_K_r10_27, u2_uk_K_r10_4, u2_uk_K_r12_15, u2_uk_K_r12_16, u2_uk_K_r3_11, u2_uk_K_r3_19, u2_uk_K_r3_4, u2_uk_K_r6_10, 
       u2_uk_K_r6_26, u2_uk_K_r6_3, u2_uk_K_r6_34, u2_uk_K_r7_13, u2_uk_K_r7_2, u2_uk_K_r7_20, u2_uk_K_r7_32, u2_uk_K_r7_39, u2_uk_K_r7_41, 
       u2_uk_K_r7_48, u2_uk_K_r7_9, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_28, u2_uk_K_r8_37, u2_uk_K_r8_42, u2_uk_K_r8_44, 
       u2_uk_K_r8_52, u2_uk_K_r8_8, u2_uk_n10, u2_uk_n100, u2_uk_n1001, u2_uk_n102, u2_uk_n1042, u2_uk_n1043, u2_uk_n1044, 
       u2_uk_n1046, u2_uk_n109, u2_uk_n11, u2_uk_n110, u2_uk_n1100, u2_uk_n1105, u2_uk_n1116, u2_uk_n1128, u2_uk_n1131, 
       u2_uk_n117, u2_uk_n118, u2_uk_n1230, u2_uk_n1236, u2_uk_n1237, u2_uk_n1245, u2_uk_n1246, u2_uk_n1251, u2_uk_n1258, 
       u2_uk_n1264, u2_uk_n1265, u2_uk_n1266, u2_uk_n1274, u2_uk_n128, u2_uk_n129, u2_uk_n1367, u2_uk_n1372, u2_uk_n1375, 
       u2_uk_n1377, u2_uk_n1378, u2_uk_n1379, u2_uk_n1381, u2_uk_n1395, u2_uk_n1396, u2_uk_n1405, u2_uk_n142, u2_uk_n145, 
       u2_uk_n146, u2_uk_n147, u2_uk_n1501, u2_uk_n1502, u2_uk_n1506, u2_uk_n1507, u2_uk_n1514, u2_uk_n1515, u2_uk_n1518, 
       u2_uk_n1519, u2_uk_n1522, u2_uk_n1529, u2_uk_n1544, u2_uk_n1568, u2_uk_n1570, u2_uk_n1573, u2_uk_n1586, u2_uk_n1594, 
       u2_uk_n1615, u2_uk_n162, u2_uk_n1622, u2_uk_n163, u2_uk_n1682, u2_uk_n1683, u2_uk_n1688, u2_uk_n1689, u2_uk_n17, 
       u2_uk_n1702, u2_uk_n1708, u2_uk_n1709, u2_uk_n1715, u2_uk_n1720, u2_uk_n1722, u2_uk_n1768, u2_uk_n1777, u2_uk_n1790, 
       u2_uk_n1799, u2_uk_n1800, u2_uk_n1802, u2_uk_n1806, u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n203, u2_uk_n207, 
       u2_uk_n222, u2_uk_n223, u2_uk_n238, u2_uk_n27, u2_uk_n299, u2_uk_n31, u2_uk_n408, u2_uk_n421, u2_uk_n500, 
       u2_uk_n520, u2_uk_n60, u2_uk_n63, u2_uk_n83, u2_uk_n93, u2_uk_n931, u2_uk_n94, u2_uk_n979, u2_uk_n984, 
       u2_uk_n986, u2_uk_n99, u0_N322, u0_N327, u0_N333, u0_N344, u0_N354, u0_N355, u0_N356, u0_N358, u0_N359, 
        u0_N362, u0_N363, u0_N365, u0_N366, u0_N370, u0_N372, u0_N373, u0_N376, u0_N378, 
        u0_N380, u0_N383, u0_N388, u0_N392, u0_N398, u0_N400, u0_N404, u0_N406, u0_N410, 
        u0_N414, u2_N0, u2_N10, u2_N11, u2_N128, u2_N129, u2_N13, u2_N130, u2_N133, 
        u2_N135, u2_N136, u2_N137, u2_N14, u2_N140, u2_N141, u2_N143, u2_N144, u2_N145, 
        u2_N147, u2_N150, u2_N151, u2_N152, u2_N153, u2_N155, u2_N157, u2_N158, u2_N18, 
        u2_N19, u2_N2, u2_N20, u2_N21, u2_N229, u2_N232, u2_N239, u2_N24, u2_N240, 
        u2_N246, u2_N247, u2_N25, u2_N253, u2_N254, u2_N256, u2_N258, u2_N26, u2_N263, 
        u2_N265, u2_N269, u2_N275, u2_N28, u2_N280, u2_N281, u2_N291, u2_N294, u2_N298, 
        u2_N299, u2_N3, u2_N306, u2_N309, u2_N31, u2_N316, u2_N319, u2_N35, u2_N353, 
        u2_N360, u2_N364, u2_N368, u2_N369, u2_N374, u2_N379, u2_N38, u2_N382, u2_N4, 
        u2_N42, u2_N420, u2_N43, u2_N430, u2_N436, u2_N442, u2_N50, u2_N53, u2_N6, 
        u2_N60, u2_N63, u2_N7, u2_N9, u2_u0_X_1, u2_uk_n1142, u2_uk_n1144, u2_uk_n1149, u2_uk_n1152, 
        u2_uk_n1167, u2_uk_n1171, u2_uk_n1178, u2_uk_n1179, u2_uk_n1183, u2_uk_n148, u2_uk_n155, u2_uk_n164, u2_uk_n182, 
        u2_uk_n202, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n231, u2_uk_n92 );
  input u0_K12_34, u0_K12_35, u0_K12_36, u0_K12_39, u0_K12_40, u0_K12_48, u0_K13_45, u0_K13_46, u0_K13_48, 
        u0_L10_11, u0_L10_12, u0_L10_14, u0_L10_15, u0_L10_19, u0_L10_21, u0_L10_22, u0_L10_25, u0_L10_27, 
        u0_L10_29, u0_L10_3, u0_L10_32, u0_L10_4, u0_L10_5, u0_L10_7, u0_L10_8, u0_L11_15, u0_L11_17, 
        u0_L11_21, u0_L11_23, u0_L11_27, u0_L11_31, u0_L11_5, u0_L11_9, u0_L9_14, u0_L9_25, u0_L9_3, 
        u0_L9_8, u0_R10_1, u0_R10_16, u0_R10_17, u0_R10_18, u0_R10_19, u0_R10_20, u0_R10_21, u0_R10_22, 
        u0_R10_23, u0_R10_24, u0_R10_25, u0_R10_26, u0_R10_27, u0_R10_28, u0_R10_29, u0_R10_30, u0_R10_31, 
        u0_R10_32, u0_R11_1, u0_R11_2, u0_R11_28, u0_R11_29, u0_R11_3, u0_R11_30, u0_R11_31, u0_R11_32, 
        u0_R11_4, u0_R11_5, u0_R9_16, u0_R9_17, u0_R9_18, u0_R9_19, u0_R9_20, u0_R9_21, u0_uk_K_r10_14, 
        u0_uk_K_r10_23, u0_uk_K_r10_28, u0_uk_K_r10_37, u0_uk_K_r10_42, u0_uk_K_r10_43, u0_uk_K_r10_44, u0_uk_K_r10_9, u0_uk_K_r11_19, u0_uk_K_r11_24, 
        u0_uk_K_r11_25, u0_uk_K_r11_26, u0_uk_K_r11_29, u0_uk_K_r11_4, u0_uk_K_r11_46, u0_uk_K_r11_48, u0_uk_K_r11_53, u0_uk_K_r9_0, u0_uk_K_r9_1, 
        u0_uk_K_r9_35, u0_uk_K_r9_9, u0_uk_n10, u0_uk_n100, u0_uk_n102, u0_uk_n106, u0_uk_n107, u0_uk_n109, u0_uk_n11, 
        u0_uk_n110, u0_uk_n117, u0_uk_n118, u0_uk_n119, u0_uk_n121, u0_uk_n126, u0_uk_n129, u0_uk_n131, u0_uk_n134, 
        u0_uk_n139, u0_uk_n140, u0_uk_n141, u0_uk_n142, u0_uk_n144, u0_uk_n145, u0_uk_n148, u0_uk_n151, u0_uk_n152, 
        u0_uk_n153, u0_uk_n154, u0_uk_n159, u0_uk_n161, u0_uk_n163, u0_uk_n167, u0_uk_n168, u0_uk_n171, u0_uk_n173, 
        u0_uk_n174, u0_uk_n178, u0_uk_n179, u0_uk_n180, u0_uk_n182, u0_uk_n184, u0_uk_n191, u0_uk_n192, u0_uk_n193, 
        u0_uk_n198, u0_uk_n203, u0_uk_n204, u0_uk_n207, u0_uk_n208, u0_uk_n211, u0_uk_n213, u0_uk_n214, u0_uk_n216, 
        u0_uk_n217, u0_uk_n220, u0_uk_n222, u0_uk_n224, u0_uk_n238, u0_uk_n242, u0_uk_n250, u0_uk_n251, u0_uk_n252, 
        u0_uk_n31, u0_uk_n60, u0_uk_n83, u0_uk_n92, u0_uk_n93, u0_uk_n94, u0_uk_n96, u0_uk_n99, u2_K10_32, 
        u2_K10_34, u2_K10_36, u2_K10_42, u2_K12_2, u2_K12_8, u2_K1_19, u2_K1_21, u2_K1_24, u2_K1_28, 
        u2_K1_37, u2_K1_40, u2_K1_43, u2_K1_45, u2_K1_46, u2_K2_34, u2_K2_35, u2_K2_36, u2_K2_40, 
        u2_K5_1, u2_K5_10, u2_K5_11, u2_K5_13, u2_K5_14, u2_K5_16, u2_K5_17, u2_K5_18, u2_K5_19, 
        u2_K5_21, u2_K5_23, u2_K5_24, u2_K5_25, u2_K5_26, u2_K5_28, u2_K5_3, u2_K5_5, u2_K5_6, 
        u2_K5_8, u2_K5_9, u2_K8_18, u2_K8_5, u2_K9_23, u2_K9_25, u2_K9_28, u2_K9_29, u2_L0_11, 
        u2_L0_12, u2_L0_19, u2_L0_22, u2_L0_29, u2_L0_32, u2_L0_4, u2_L0_7, u2_L10_13, u2_L10_17, 
        u2_L10_18, u2_L10_2, u2_L10_23, u2_L10_28, u2_L10_31, u2_L10_9, u2_L12_15, u2_L12_21, u2_L12_27, 
        u2_L12_5, u2_L3_1, u2_L3_10, u2_L3_13, u2_L3_14, u2_L3_16, u2_L3_17, u2_L3_18, u2_L3_2, 
        u2_L3_20, u2_L3_23, u2_L3_24, u2_L3_25, u2_L3_26, u2_L3_28, u2_L3_3, u2_L3_30, u2_L3_31, 
        u2_L3_6, u2_L3_8, u2_L3_9, u2_L6_16, u2_L6_17, u2_L6_23, u2_L6_24, u2_L6_30, u2_L6_31, 
        u2_L6_6, u2_L6_9, u2_L7_1, u2_L7_10, u2_L7_14, u2_L7_20, u2_L7_25, u2_L7_26, u2_L7_3, 
        u2_L7_8, u2_L8_11, u2_L8_12, u2_L8_19, u2_L8_22, u2_L8_29, u2_L8_32, u2_L8_4, u2_L8_7, 
        u2_R0_20, u2_R0_21, u2_R0_22, u2_R0_23, u2_R0_24, u2_R0_25, u2_R0_26, u2_R0_27, u2_R0_28, 
        u2_R0_29, u2_R10_1, u2_R10_2, u2_R10_3, u2_R10_32, u2_R10_4, u2_R10_5, u2_R10_6, u2_R10_7, 
        u2_R10_8, u2_R10_9, u2_R12_1, u2_R12_28, u2_R12_29, u2_R12_30, u2_R12_31, u2_R12_32, u2_R3_1, 
        u2_R3_10, u2_R3_11, u2_R3_12, u2_R3_13, u2_R3_14, u2_R3_15, u2_R3_16, u2_R3_17, u2_R3_18, 
        u2_R3_19, u2_R3_2, u2_R3_20, u2_R3_21, u2_R3_3, u2_R3_32, u2_R3_4, u2_R3_5, u2_R3_6, 
        u2_R3_7, u2_R3_8, u2_R3_9, u2_R6_1, u2_R6_10, u2_R6_11, u2_R6_12, u2_R6_13, u2_R6_2, 
        u2_R6_3, u2_R6_32, u2_R6_4, u2_R6_5, u2_R6_8, u2_R6_9, u2_R7_12, u2_R7_13, u2_R7_14, 
        u2_R7_15, u2_R7_16, u2_R7_17, u2_R7_18, u2_R7_19, u2_R7_20, u2_R7_21, u2_R8_20, u2_R8_21, 
        u2_R8_22, u2_R8_23, u2_R8_24, u2_R8_25, u2_R8_26, u2_R8_27, u2_R8_28, u2_R8_29, u2_desIn_r_0, 
        u2_desIn_r_1, u2_desIn_r_11, u2_desIn_r_12, u2_desIn_r_16, u2_desIn_r_17, u2_desIn_r_18, u2_desIn_r_19, u2_desIn_r_20, u2_desIn_r_22, 
        u2_desIn_r_25, u2_desIn_r_26, u2_desIn_r_27, u2_desIn_r_28, u2_desIn_r_29, u2_desIn_r_3, u2_desIn_r_30, u2_desIn_r_32, u2_desIn_r_33, 
        u2_desIn_r_34, u2_desIn_r_35, u2_desIn_r_37, u2_desIn_r_38, u2_desIn_r_41, u2_desIn_r_42, u2_desIn_r_43, u2_desIn_r_44, u2_desIn_r_45, 
        u2_desIn_r_49, u2_desIn_r_51, u2_desIn_r_52, u2_desIn_r_53, u2_desIn_r_54, u2_desIn_r_56, u2_desIn_r_57, u2_desIn_r_59, u2_desIn_r_6, 
        u2_desIn_r_61, u2_desIn_r_62, u2_desIn_r_7, u2_desIn_r_8, u2_desIn_r_9, u2_key_r_0, u2_key_r_14, u2_key_r_16, u2_key_r_2, 
        u2_key_r_21, u2_key_r_22, u2_key_r_23, u2_key_r_25, u2_key_r_28, u2_key_r_29, u2_key_r_30, u2_key_r_31, u2_key_r_32, 
        u2_key_r_33, u2_key_r_35, u2_key_r_36, u2_key_r_37, u2_key_r_40, u2_key_r_42, u2_key_r_43, u2_key_r_44, u2_key_r_47, 
        u2_key_r_48, u2_key_r_51, u2_key_r_52, u2_key_r_55, u2_key_r_7, u2_key_r_9, u2_uk_K_r0_15, u2_uk_K_r0_31, u2_uk_K_r0_36, 
        u2_uk_K_r10_10, u2_uk_K_r10_27, u2_uk_K_r10_4, u2_uk_K_r12_15, u2_uk_K_r12_16, u2_uk_K_r3_11, u2_uk_K_r3_19, u2_uk_K_r3_4, u2_uk_K_r6_10, 
        u2_uk_K_r6_26, u2_uk_K_r6_3, u2_uk_K_r6_34, u2_uk_K_r7_13, u2_uk_K_r7_2, u2_uk_K_r7_20, u2_uk_K_r7_32, u2_uk_K_r7_39, u2_uk_K_r7_41, 
        u2_uk_K_r7_48, u2_uk_K_r7_9, u2_uk_K_r8_16, u2_uk_K_r8_2, u2_uk_K_r8_22, u2_uk_K_r8_28, u2_uk_K_r8_37, u2_uk_K_r8_42, u2_uk_K_r8_44, 
        u2_uk_K_r8_52, u2_uk_K_r8_8, u2_uk_n10, u2_uk_n100, u2_uk_n1001, u2_uk_n102, u2_uk_n1042, u2_uk_n1043, u2_uk_n1044, 
        u2_uk_n1046, u2_uk_n109, u2_uk_n11, u2_uk_n110, u2_uk_n1100, u2_uk_n1105, u2_uk_n1116, u2_uk_n1128, u2_uk_n1131, 
        u2_uk_n117, u2_uk_n118, u2_uk_n1230, u2_uk_n1236, u2_uk_n1237, u2_uk_n1245, u2_uk_n1246, u2_uk_n1251, u2_uk_n1258, 
        u2_uk_n1264, u2_uk_n1265, u2_uk_n1266, u2_uk_n1274, u2_uk_n128, u2_uk_n129, u2_uk_n1367, u2_uk_n1372, u2_uk_n1375, 
        u2_uk_n1377, u2_uk_n1378, u2_uk_n1379, u2_uk_n1381, u2_uk_n1395, u2_uk_n1396, u2_uk_n1405, u2_uk_n142, u2_uk_n145, 
        u2_uk_n146, u2_uk_n147, u2_uk_n1501, u2_uk_n1502, u2_uk_n1506, u2_uk_n1507, u2_uk_n1514, u2_uk_n1515, u2_uk_n1518, 
        u2_uk_n1519, u2_uk_n1522, u2_uk_n1529, u2_uk_n1544, u2_uk_n1568, u2_uk_n1570, u2_uk_n1573, u2_uk_n1586, u2_uk_n1594, 
        u2_uk_n1615, u2_uk_n162, u2_uk_n1622, u2_uk_n163, u2_uk_n1682, u2_uk_n1683, u2_uk_n1688, u2_uk_n1689, u2_uk_n17, 
        u2_uk_n1702, u2_uk_n1708, u2_uk_n1709, u2_uk_n1715, u2_uk_n1720, u2_uk_n1722, u2_uk_n1768, u2_uk_n1777, u2_uk_n1790, 
        u2_uk_n1799, u2_uk_n1800, u2_uk_n1802, u2_uk_n1806, u2_uk_n187, u2_uk_n188, u2_uk_n191, u2_uk_n203, u2_uk_n207, 
        u2_uk_n222, u2_uk_n223, u2_uk_n238, u2_uk_n27, u2_uk_n299, u2_uk_n31, u2_uk_n408, u2_uk_n421, u2_uk_n500, 
        u2_uk_n520, u2_uk_n60, u2_uk_n63, u2_uk_n83, u2_uk_n93, u2_uk_n931, u2_uk_n94, u2_uk_n979, u2_uk_n984, 
        u2_uk_n986, u2_uk_n99;
  output u0_N322, u0_N327, u0_N333, u0_N344, u0_N354, u0_N355, u0_N356, u0_N358, u0_N359, 
        u0_N362, u0_N363, u0_N365, u0_N366, u0_N370, u0_N372, u0_N373, u0_N376, u0_N378, 
        u0_N380, u0_N383, u0_N388, u0_N392, u0_N398, u0_N400, u0_N404, u0_N406, u0_N410, 
        u0_N414, u2_N0, u2_N10, u2_N11, u2_N128, u2_N129, u2_N13, u2_N130, u2_N133, 
        u2_N135, u2_N136, u2_N137, u2_N14, u2_N140, u2_N141, u2_N143, u2_N144, u2_N145, 
        u2_N147, u2_N150, u2_N151, u2_N152, u2_N153, u2_N155, u2_N157, u2_N158, u2_N18, 
        u2_N19, u2_N2, u2_N20, u2_N21, u2_N229, u2_N232, u2_N239, u2_N24, u2_N240, 
        u2_N246, u2_N247, u2_N25, u2_N253, u2_N254, u2_N256, u2_N258, u2_N26, u2_N263, 
        u2_N265, u2_N269, u2_N275, u2_N28, u2_N280, u2_N281, u2_N291, u2_N294, u2_N298, 
        u2_N299, u2_N3, u2_N306, u2_N309, u2_N31, u2_N316, u2_N319, u2_N35, u2_N353, 
        u2_N360, u2_N364, u2_N368, u2_N369, u2_N374, u2_N379, u2_N38, u2_N382, u2_N4, 
        u2_N42, u2_N420, u2_N43, u2_N430, u2_N436, u2_N442, u2_N50, u2_N53, u2_N6, 
        u2_N60, u2_N63, u2_N7, u2_N9, u2_u0_X_1, u2_uk_n1142, u2_uk_n1144, u2_uk_n1149, u2_uk_n1152, 
        u2_uk_n1167, u2_uk_n1171, u2_uk_n1178, u2_uk_n1179, u2_uk_n1183, u2_uk_n148, u2_uk_n155, u2_uk_n164, u2_uk_n182, 
        u2_uk_n202, u2_uk_n208, u2_uk_n209, u2_uk_n213, u2_uk_n214, u2_uk_n217, u2_uk_n220, u2_uk_n231, u2_uk_n92;
  wire u0_K11_25, u0_K11_26, u0_K11_27, u0_K11_28, u0_K11_29, u0_K11_30, u0_K12_25, u0_K12_26, u0_K12_27, 
       u0_K12_28, u0_K12_29, u0_K12_30, u0_K12_31, u0_K12_32, u0_K12_33, u0_K12_37, u0_K12_38, u0_K12_41, 
       u0_K12_42, u0_K12_43, u0_K12_44, u0_K12_45, u0_K12_46, u0_K12_47, u0_K13_1, u0_K13_2, u0_K13_3, 
       u0_K13_4, u0_K13_43, u0_K13_44, u0_K13_47, u0_K13_5, u0_K13_6, u0_out10_14, u0_out10_25, u0_out10_3, 
       u0_out10_8, u0_out11_11, u0_out11_12, u0_out11_14, u0_out11_15, u0_out11_19, u0_out11_21, u0_out11_22, u0_out11_25, 
       u0_out11_27, u0_out11_29, u0_out11_3, u0_out11_32, u0_out11_4, u0_out11_5, u0_out11_7, u0_out11_8, u0_out12_15, 
       u0_out12_17, u0_out12_21, u0_out12_23, u0_out12_27, u0_out12_31, u0_out12_5, u0_out12_9, u0_u10_X_25, u0_u10_X_26, 
       u0_u10_X_27, u0_u10_X_28, u0_u10_X_29, u0_u10_X_30, u0_u10_u4_n100, u0_u10_u4_n101, u0_u10_u4_n102, u0_u10_u4_n103, u0_u10_u4_n104, 
       u0_u10_u4_n105, u0_u10_u4_n106, u0_u10_u4_n107, u0_u10_u4_n108, u0_u10_u4_n109, u0_u10_u4_n110, u0_u10_u4_n111, u0_u10_u4_n112, u0_u10_u4_n113, 
       u0_u10_u4_n114, u0_u10_u4_n115, u0_u10_u4_n116, u0_u10_u4_n117, u0_u10_u4_n118, u0_u10_u4_n119, u0_u10_u4_n120, u0_u10_u4_n121, u0_u10_u4_n122, 
       u0_u10_u4_n123, u0_u10_u4_n124, u0_u10_u4_n125, u0_u10_u4_n126, u0_u10_u4_n127, u0_u10_u4_n128, u0_u10_u4_n129, u0_u10_u4_n130, u0_u10_u4_n131, 
       u0_u10_u4_n132, u0_u10_u4_n133, u0_u10_u4_n134, u0_u10_u4_n135, u0_u10_u4_n136, u0_u10_u4_n137, u0_u10_u4_n138, u0_u10_u4_n139, u0_u10_u4_n140, 
       u0_u10_u4_n141, u0_u10_u4_n142, u0_u10_u4_n143, u0_u10_u4_n144, u0_u10_u4_n145, u0_u10_u4_n146, u0_u10_u4_n147, u0_u10_u4_n148, u0_u10_u4_n149, 
       u0_u10_u4_n150, u0_u10_u4_n151, u0_u10_u4_n152, u0_u10_u4_n153, u0_u10_u4_n154, u0_u10_u4_n155, u0_u10_u4_n156, u0_u10_u4_n157, u0_u10_u4_n158, 
       u0_u10_u4_n159, u0_u10_u4_n160, u0_u10_u4_n161, u0_u10_u4_n162, u0_u10_u4_n163, u0_u10_u4_n164, u0_u10_u4_n165, u0_u10_u4_n166, u0_u10_u4_n167, 
       u0_u10_u4_n168, u0_u10_u4_n169, u0_u10_u4_n170, u0_u10_u4_n171, u0_u10_u4_n172, u0_u10_u4_n173, u0_u10_u4_n174, u0_u10_u4_n175, u0_u10_u4_n176, 
       u0_u10_u4_n177, u0_u10_u4_n178, u0_u10_u4_n179, u0_u10_u4_n180, u0_u10_u4_n181, u0_u10_u4_n182, u0_u10_u4_n183, u0_u10_u4_n184, u0_u10_u4_n185, 
       u0_u10_u4_n186, u0_u10_u4_n94, u0_u10_u4_n95, u0_u10_u4_n96, u0_u10_u4_n97, u0_u10_u4_n98, u0_u10_u4_n99, u0_u11_X_25, u0_u11_X_26, 
       u0_u11_X_27, u0_u11_X_28, u0_u11_X_29, u0_u11_X_30, u0_u11_X_31, u0_u11_X_32, u0_u11_X_33, u0_u11_X_34, u0_u11_X_35, 
       u0_u11_X_36, u0_u11_X_37, u0_u11_X_38, u0_u11_X_39, u0_u11_X_40, u0_u11_X_41, u0_u11_X_42, u0_u11_X_43, u0_u11_X_44, 
       u0_u11_X_45, u0_u11_X_46, u0_u11_X_47, u0_u11_X_48, u0_u11_u4_n100, u0_u11_u4_n101, u0_u11_u4_n102, u0_u11_u4_n103, u0_u11_u4_n104, 
       u0_u11_u4_n105, u0_u11_u4_n106, u0_u11_u4_n107, u0_u11_u4_n108, u0_u11_u4_n109, u0_u11_u4_n110, u0_u11_u4_n111, u0_u11_u4_n112, u0_u11_u4_n113, 
       u0_u11_u4_n114, u0_u11_u4_n115, u0_u11_u4_n116, u0_u11_u4_n117, u0_u11_u4_n118, u0_u11_u4_n119, u0_u11_u4_n120, u0_u11_u4_n121, u0_u11_u4_n122, 
       u0_u11_u4_n123, u0_u11_u4_n124, u0_u11_u4_n125, u0_u11_u4_n126, u0_u11_u4_n127, u0_u11_u4_n128, u0_u11_u4_n129, u0_u11_u4_n130, u0_u11_u4_n131, 
       u0_u11_u4_n132, u0_u11_u4_n133, u0_u11_u4_n134, u0_u11_u4_n135, u0_u11_u4_n136, u0_u11_u4_n137, u0_u11_u4_n138, u0_u11_u4_n139, u0_u11_u4_n140, 
       u0_u11_u4_n141, u0_u11_u4_n142, u0_u11_u4_n143, u0_u11_u4_n144, u0_u11_u4_n145, u0_u11_u4_n146, u0_u11_u4_n147, u0_u11_u4_n148, u0_u11_u4_n149, 
       u0_u11_u4_n150, u0_u11_u4_n151, u0_u11_u4_n152, u0_u11_u4_n153, u0_u11_u4_n154, u0_u11_u4_n155, u0_u11_u4_n156, u0_u11_u4_n157, u0_u11_u4_n158, 
       u0_u11_u4_n159, u0_u11_u4_n160, u0_u11_u4_n161, u0_u11_u4_n162, u0_u11_u4_n163, u0_u11_u4_n164, u0_u11_u4_n165, u0_u11_u4_n166, u0_u11_u4_n167, 
       u0_u11_u4_n168, u0_u11_u4_n169, u0_u11_u4_n170, u0_u11_u4_n171, u0_u11_u4_n172, u0_u11_u4_n173, u0_u11_u4_n174, u0_u11_u4_n175, u0_u11_u4_n176, 
       u0_u11_u4_n177, u0_u11_u4_n178, u0_u11_u4_n179, u0_u11_u4_n180, u0_u11_u4_n181, u0_u11_u4_n182, u0_u11_u4_n183, u0_u11_u4_n184, u0_u11_u4_n185, 
       u0_u11_u4_n186, u0_u11_u4_n94, u0_u11_u4_n95, u0_u11_u4_n96, u0_u11_u4_n97, u0_u11_u4_n98, u0_u11_u4_n99, u0_u11_u5_n100, u0_u11_u5_n101, 
       u0_u11_u5_n102, u0_u11_u5_n103, u0_u11_u5_n104, u0_u11_u5_n105, u0_u11_u5_n106, u0_u11_u5_n107, u0_u11_u5_n108, u0_u11_u5_n109, u0_u11_u5_n110, 
       u0_u11_u5_n111, u0_u11_u5_n112, u0_u11_u5_n113, u0_u11_u5_n114, u0_u11_u5_n115, u0_u11_u5_n116, u0_u11_u5_n117, u0_u11_u5_n118, u0_u11_u5_n119, 
       u0_u11_u5_n120, u0_u11_u5_n121, u0_u11_u5_n122, u0_u11_u5_n123, u0_u11_u5_n124, u0_u11_u5_n125, u0_u11_u5_n126, u0_u11_u5_n127, u0_u11_u5_n128, 
       u0_u11_u5_n129, u0_u11_u5_n130, u0_u11_u5_n131, u0_u11_u5_n132, u0_u11_u5_n133, u0_u11_u5_n134, u0_u11_u5_n135, u0_u11_u5_n136, u0_u11_u5_n137, 
       u0_u11_u5_n138, u0_u11_u5_n139, u0_u11_u5_n140, u0_u11_u5_n141, u0_u11_u5_n142, u0_u11_u5_n143, u0_u11_u5_n144, u0_u11_u5_n145, u0_u11_u5_n146, 
       u0_u11_u5_n147, u0_u11_u5_n148, u0_u11_u5_n149, u0_u11_u5_n150, u0_u11_u5_n151, u0_u11_u5_n152, u0_u11_u5_n153, u0_u11_u5_n154, u0_u11_u5_n155, 
       u0_u11_u5_n156, u0_u11_u5_n157, u0_u11_u5_n158, u0_u11_u5_n159, u0_u11_u5_n160, u0_u11_u5_n161, u0_u11_u5_n162, u0_u11_u5_n163, u0_u11_u5_n164, 
       u0_u11_u5_n165, u0_u11_u5_n166, u0_u11_u5_n167, u0_u11_u5_n168, u0_u11_u5_n169, u0_u11_u5_n170, u0_u11_u5_n171, u0_u11_u5_n172, u0_u11_u5_n173, 
       u0_u11_u5_n174, u0_u11_u5_n175, u0_u11_u5_n176, u0_u11_u5_n177, u0_u11_u5_n178, u0_u11_u5_n179, u0_u11_u5_n180, u0_u11_u5_n181, u0_u11_u5_n182, 
       u0_u11_u5_n183, u0_u11_u5_n184, u0_u11_u5_n185, u0_u11_u5_n186, u0_u11_u5_n187, u0_u11_u5_n188, u0_u11_u5_n189, u0_u11_u5_n190, u0_u11_u5_n191, 
       u0_u11_u5_n192, u0_u11_u5_n193, u0_u11_u5_n194, u0_u11_u5_n195, u0_u11_u5_n196, u0_u11_u5_n99, u0_u11_u6_n100, u0_u11_u6_n101, u0_u11_u6_n102, 
       u0_u11_u6_n103, u0_u11_u6_n104, u0_u11_u6_n105, u0_u11_u6_n106, u0_u11_u6_n107, u0_u11_u6_n108, u0_u11_u6_n109, u0_u11_u6_n110, u0_u11_u6_n111, 
       u0_u11_u6_n112, u0_u11_u6_n113, u0_u11_u6_n114, u0_u11_u6_n115, u0_u11_u6_n116, u0_u11_u6_n117, u0_u11_u6_n118, u0_u11_u6_n119, u0_u11_u6_n120, 
       u0_u11_u6_n121, u0_u11_u6_n122, u0_u11_u6_n123, u0_u11_u6_n124, u0_u11_u6_n125, u0_u11_u6_n126, u0_u11_u6_n127, u0_u11_u6_n128, u0_u11_u6_n129, 
       u0_u11_u6_n130, u0_u11_u6_n131, u0_u11_u6_n132, u0_u11_u6_n133, u0_u11_u6_n134, u0_u11_u6_n135, u0_u11_u6_n136, u0_u11_u6_n137, u0_u11_u6_n138, 
       u0_u11_u6_n139, u0_u11_u6_n140, u0_u11_u6_n141, u0_u11_u6_n142, u0_u11_u6_n143, u0_u11_u6_n144, u0_u11_u6_n145, u0_u11_u6_n146, u0_u11_u6_n147, 
       u0_u11_u6_n148, u0_u11_u6_n149, u0_u11_u6_n150, u0_u11_u6_n151, u0_u11_u6_n152, u0_u11_u6_n153, u0_u11_u6_n154, u0_u11_u6_n155, u0_u11_u6_n156, 
       u0_u11_u6_n157, u0_u11_u6_n158, u0_u11_u6_n159, u0_u11_u6_n160, u0_u11_u6_n161, u0_u11_u6_n162, u0_u11_u6_n163, u0_u11_u6_n164, u0_u11_u6_n165, 
       u0_u11_u6_n166, u0_u11_u6_n167, u0_u11_u6_n168, u0_u11_u6_n169, u0_u11_u6_n170, u0_u11_u6_n171, u0_u11_u6_n172, u0_u11_u6_n173, u0_u11_u6_n174, 
       u0_u11_u6_n88, u0_u11_u6_n89, u0_u11_u6_n90, u0_u11_u6_n91, u0_u11_u6_n92, u0_u11_u6_n93, u0_u11_u6_n94, u0_u11_u6_n95, u0_u11_u6_n96, 
       u0_u11_u6_n97, u0_u11_u6_n98, u0_u11_u6_n99, u0_u11_u7_n100, u0_u11_u7_n101, u0_u11_u7_n102, u0_u11_u7_n103, u0_u11_u7_n104, u0_u11_u7_n105, 
       u0_u11_u7_n106, u0_u11_u7_n107, u0_u11_u7_n108, u0_u11_u7_n109, u0_u11_u7_n110, u0_u11_u7_n111, u0_u11_u7_n112, u0_u11_u7_n113, u0_u11_u7_n114, 
       u0_u11_u7_n115, u0_u11_u7_n116, u0_u11_u7_n117, u0_u11_u7_n118, u0_u11_u7_n119, u0_u11_u7_n120, u0_u11_u7_n121, u0_u11_u7_n122, u0_u11_u7_n123, 
       u0_u11_u7_n124, u0_u11_u7_n125, u0_u11_u7_n126, u0_u11_u7_n127, u0_u11_u7_n128, u0_u11_u7_n129, u0_u11_u7_n130, u0_u11_u7_n131, u0_u11_u7_n132, 
       u0_u11_u7_n133, u0_u11_u7_n134, u0_u11_u7_n135, u0_u11_u7_n136, u0_u11_u7_n137, u0_u11_u7_n138, u0_u11_u7_n139, u0_u11_u7_n140, u0_u11_u7_n141, 
       u0_u11_u7_n142, u0_u11_u7_n143, u0_u11_u7_n144, u0_u11_u7_n145, u0_u11_u7_n146, u0_u11_u7_n147, u0_u11_u7_n148, u0_u11_u7_n149, u0_u11_u7_n150, 
       u0_u11_u7_n151, u0_u11_u7_n152, u0_u11_u7_n153, u0_u11_u7_n154, u0_u11_u7_n155, u0_u11_u7_n156, u0_u11_u7_n157, u0_u11_u7_n158, u0_u11_u7_n159, 
       u0_u11_u7_n160, u0_u11_u7_n161, u0_u11_u7_n162, u0_u11_u7_n163, u0_u11_u7_n164, u0_u11_u7_n165, u0_u11_u7_n166, u0_u11_u7_n167, u0_u11_u7_n168, 
       u0_u11_u7_n169, u0_u11_u7_n170, u0_u11_u7_n171, u0_u11_u7_n172, u0_u11_u7_n173, u0_u11_u7_n174, u0_u11_u7_n175, u0_u11_u7_n176, u0_u11_u7_n177, 
       u0_u11_u7_n178, u0_u11_u7_n179, u0_u11_u7_n180, u0_u11_u7_n91, u0_u11_u7_n92, u0_u11_u7_n93, u0_u11_u7_n94, u0_u11_u7_n95, u0_u11_u7_n96, 
       u0_u11_u7_n97, u0_u11_u7_n98, u0_u11_u7_n99, u0_u12_X_1, u0_u12_X_2, u0_u12_X_3, u0_u12_X_4, u0_u12_X_43, u0_u12_X_44, 
       u0_u12_X_45, u0_u12_X_46, u0_u12_X_47, u0_u12_X_48, u0_u12_X_5, u0_u12_X_6, u0_u12_u0_n100, u0_u12_u0_n101, u0_u12_u0_n102, 
       u0_u12_u0_n103, u0_u12_u0_n104, u0_u12_u0_n105, u0_u12_u0_n106, u0_u12_u0_n107, u0_u12_u0_n108, u0_u12_u0_n109, u0_u12_u0_n110, u0_u12_u0_n111, 
       u0_u12_u0_n112, u0_u12_u0_n113, u0_u12_u0_n114, u0_u12_u0_n115, u0_u12_u0_n116, u0_u12_u0_n117, u0_u12_u0_n118, u0_u12_u0_n119, u0_u12_u0_n120, 
       u0_u12_u0_n121, u0_u12_u0_n122, u0_u12_u0_n123, u0_u12_u0_n124, u0_u12_u0_n125, u0_u12_u0_n126, u0_u12_u0_n127, u0_u12_u0_n128, u0_u12_u0_n129, 
       u0_u12_u0_n130, u0_u12_u0_n131, u0_u12_u0_n132, u0_u12_u0_n133, u0_u12_u0_n134, u0_u12_u0_n135, u0_u12_u0_n136, u0_u12_u0_n137, u0_u12_u0_n138, 
       u0_u12_u0_n139, u0_u12_u0_n140, u0_u12_u0_n141, u0_u12_u0_n142, u0_u12_u0_n143, u0_u12_u0_n144, u0_u12_u0_n145, u0_u12_u0_n146, u0_u12_u0_n147, 
       u0_u12_u0_n148, u0_u12_u0_n149, u0_u12_u0_n150, u0_u12_u0_n151, u0_u12_u0_n152, u0_u12_u0_n153, u0_u12_u0_n154, u0_u12_u0_n155, u0_u12_u0_n156, 
       u0_u12_u0_n157, u0_u12_u0_n158, u0_u12_u0_n159, u0_u12_u0_n160, u0_u12_u0_n161, u0_u12_u0_n162, u0_u12_u0_n163, u0_u12_u0_n164, u0_u12_u0_n165, 
       u0_u12_u0_n166, u0_u12_u0_n167, u0_u12_u0_n168, u0_u12_u0_n169, u0_u12_u0_n170, u0_u12_u0_n171, u0_u12_u0_n172, u0_u12_u0_n173, u0_u12_u0_n174, 
       u0_u12_u0_n88, u0_u12_u0_n89, u0_u12_u0_n90, u0_u12_u0_n91, u0_u12_u0_n92, u0_u12_u0_n93, u0_u12_u0_n94, u0_u12_u0_n95, u0_u12_u0_n96, 
       u0_u12_u0_n97, u0_u12_u0_n98, u0_u12_u0_n99, u0_u12_u7_n100, u0_u12_u7_n101, u0_u12_u7_n102, u0_u12_u7_n103, u0_u12_u7_n104, u0_u12_u7_n105, 
       u0_u12_u7_n106, u0_u12_u7_n107, u0_u12_u7_n108, u0_u12_u7_n109, u0_u12_u7_n110, u0_u12_u7_n111, u0_u12_u7_n112, u0_u12_u7_n113, u0_u12_u7_n114, 
       u0_u12_u7_n115, u0_u12_u7_n116, u0_u12_u7_n117, u0_u12_u7_n118, u0_u12_u7_n119, u0_u12_u7_n120, u0_u12_u7_n121, u0_u12_u7_n122, u0_u12_u7_n123, 
       u0_u12_u7_n124, u0_u12_u7_n125, u0_u12_u7_n126, u0_u12_u7_n127, u0_u12_u7_n128, u0_u12_u7_n129, u0_u12_u7_n130, u0_u12_u7_n131, u0_u12_u7_n132, 
       u0_u12_u7_n133, u0_u12_u7_n134, u0_u12_u7_n135, u0_u12_u7_n136, u0_u12_u7_n137, u0_u12_u7_n138, u0_u12_u7_n139, u0_u12_u7_n140, u0_u12_u7_n141, 
       u0_u12_u7_n142, u0_u12_u7_n143, u0_u12_u7_n144, u0_u12_u7_n145, u0_u12_u7_n146, u0_u12_u7_n147, u0_u12_u7_n148, u0_u12_u7_n149, u0_u12_u7_n150, 
       u0_u12_u7_n151, u0_u12_u7_n152, u0_u12_u7_n153, u0_u12_u7_n154, u0_u12_u7_n155, u0_u12_u7_n156, u0_u12_u7_n157, u0_u12_u7_n158, u0_u12_u7_n159, 
       u0_u12_u7_n160, u0_u12_u7_n161, u0_u12_u7_n162, u0_u12_u7_n163, u0_u12_u7_n164, u0_u12_u7_n165, u0_u12_u7_n166, u0_u12_u7_n167, u0_u12_u7_n168, 
       u0_u12_u7_n169, u0_u12_u7_n170, u0_u12_u7_n171, u0_u12_u7_n172, u0_u12_u7_n173, u0_u12_u7_n174, u0_u12_u7_n175, u0_u12_u7_n176, u0_u12_u7_n177, 
       u0_u12_u7_n178, u0_u12_u7_n179, u0_u12_u7_n180, u0_u12_u7_n91, u0_u12_u7_n92, u0_u12_u7_n93, u0_u12_u7_n94, u0_u12_u7_n95, u0_u12_u7_n96, 
       u0_u12_u7_n97, u0_u12_u7_n98, u0_u12_u7_n99, u0_uk_n940, u0_uk_n941, u0_uk_n943, u0_uk_n944, u0_uk_n946, u0_uk_n952, 
       u0_uk_n964, u0_uk_n965, u0_uk_n966, u0_uk_n971, u0_uk_n972, u0_uk_n973, u0_uk_n974, u0_uk_n993, u0_uk_n994, 
       u0_uk_n995, u2_K10_31, u2_K10_33, u2_K10_35, u2_K10_37, u2_K10_38, u2_K10_39, u2_K10_40, u2_K10_41, 
       u2_K12_1, u2_K12_10, u2_K12_11, u2_K12_12, u2_K12_3, u2_K12_4, u2_K12_5, u2_K12_6, u2_K12_7, 
       u2_K12_9, u2_K14_43, u2_K14_44, u2_K14_45, u2_K14_46, u2_K14_47, u2_K14_48, u2_K1_1, u2_K1_20, 
       u2_K1_22, u2_K1_23, u2_K1_25, u2_K1_26, u2_K1_27, u2_K1_29, u2_K1_30, u2_K1_31, u2_K1_32, 
       u2_K1_33, u2_K1_34, u2_K1_35, u2_K1_36, u2_K1_38, u2_K1_39, u2_K1_41, u2_K1_42, u2_K1_44, 
       u2_K1_47, u2_K1_48, u2_K2_31, u2_K2_32, u2_K2_33, u2_K2_37, u2_K2_38, u2_K2_39, u2_K2_41, 
       u2_K2_42, u2_K5_12, u2_K5_15, u2_K5_2, u2_K5_20, u2_K5_22, u2_K5_27, u2_K5_29, u2_K5_30, 
       u2_K5_4, u2_K5_7, u2_K8_1, u2_K8_13, u2_K8_14, u2_K8_15, u2_K8_16, u2_K8_17, u2_K8_2, 
       u2_K8_3, u2_K8_4, u2_K8_6, u2_K9_19, u2_K9_20, u2_K9_21, u2_K9_22, u2_K9_24, u2_K9_26, 
       u2_K9_27, u2_K9_30, u2_out0_1, u2_out0_10, u2_out0_11, u2_out0_12, u2_out0_14, u2_out0_15, u2_out0_19, 
       u2_out0_20, u2_out0_21, u2_out0_22, u2_out0_25, u2_out0_26, u2_out0_27, u2_out0_29, u2_out0_3, u2_out0_32, 
       u2_out0_4, u2_out0_5, u2_out0_7, u2_out0_8, u2_out11_13, u2_out11_17, u2_out11_18, u2_out11_2, u2_out11_23, 
       u2_out11_28, u2_out11_31, u2_out11_9, u2_out13_15, u2_out13_21, u2_out13_27, u2_out13_5, u2_out1_11, u2_out1_12, 
       u2_out1_19, u2_out1_22, u2_out1_29, u2_out1_32, u2_out1_4, u2_out1_7, u2_out4_1, u2_out4_10, u2_out4_13, 
       u2_out4_14, u2_out4_16, u2_out4_17, u2_out4_18, u2_out4_2, u2_out4_20, u2_out4_23, u2_out4_24, u2_out4_25, 
       u2_out4_26, u2_out4_28, u2_out4_3, u2_out4_30, u2_out4_31, u2_out4_6, u2_out4_8, u2_out4_9, u2_out7_16, 
       u2_out7_17, u2_out7_23, u2_out7_24, u2_out7_30, u2_out7_31, u2_out7_6, u2_out7_9, u2_out8_1, u2_out8_10, 
       u2_out8_14, u2_out8_20, u2_out8_25, u2_out8_26, u2_out8_3, u2_out8_8, u2_out9_11, u2_out9_12, u2_out9_19, 
       u2_out9_22, u2_out9_29, u2_out9_32, u2_out9_4, u2_out9_7, u2_u0_X_19, u2_u0_X_20, u2_u0_X_21, u2_u0_X_22, 
       u2_u0_X_23, u2_u0_X_24, u2_u0_X_25, u2_u0_X_26, u2_u0_X_27, u2_u0_X_28, u2_u0_X_29, u2_u0_X_30, u2_u0_X_31, 
       u2_u0_X_32, u2_u0_X_33, u2_u0_X_34, u2_u0_X_35, u2_u0_X_36, u2_u0_X_37, u2_u0_X_38, u2_u0_X_39, u2_u0_X_40, 
       u2_u0_X_41, u2_u0_X_42, u2_u0_X_43, u2_u0_X_44, u2_u0_X_45, u2_u0_X_46, u2_u0_X_47, u2_u0_X_48, u2_u0_u3_n100, 
       u2_u0_u3_n101, u2_u0_u3_n102, u2_u0_u3_n103, u2_u0_u3_n104, u2_u0_u3_n105, u2_u0_u3_n106, u2_u0_u3_n107, u2_u0_u3_n108, u2_u0_u3_n109, 
       u2_u0_u3_n110, u2_u0_u3_n111, u2_u0_u3_n112, u2_u0_u3_n113, u2_u0_u3_n114, u2_u0_u3_n115, u2_u0_u3_n116, u2_u0_u3_n117, u2_u0_u3_n118, 
       u2_u0_u3_n119, u2_u0_u3_n120, u2_u0_u3_n121, u2_u0_u3_n122, u2_u0_u3_n123, u2_u0_u3_n124, u2_u0_u3_n125, u2_u0_u3_n126, u2_u0_u3_n127, 
       u2_u0_u3_n128, u2_u0_u3_n129, u2_u0_u3_n130, u2_u0_u3_n131, u2_u0_u3_n132, u2_u0_u3_n133, u2_u0_u3_n134, u2_u0_u3_n135, u2_u0_u3_n136, 
       u2_u0_u3_n137, u2_u0_u3_n138, u2_u0_u3_n139, u2_u0_u3_n140, u2_u0_u3_n141, u2_u0_u3_n142, u2_u0_u3_n143, u2_u0_u3_n144, u2_u0_u3_n145, 
       u2_u0_u3_n146, u2_u0_u3_n147, u2_u0_u3_n148, u2_u0_u3_n149, u2_u0_u3_n150, u2_u0_u3_n151, u2_u0_u3_n152, u2_u0_u3_n153, u2_u0_u3_n154, 
       u2_u0_u3_n155, u2_u0_u3_n156, u2_u0_u3_n157, u2_u0_u3_n158, u2_u0_u3_n159, u2_u0_u3_n160, u2_u0_u3_n161, u2_u0_u3_n162, u2_u0_u3_n163, 
       u2_u0_u3_n164, u2_u0_u3_n165, u2_u0_u3_n166, u2_u0_u3_n167, u2_u0_u3_n168, u2_u0_u3_n169, u2_u0_u3_n170, u2_u0_u3_n171, u2_u0_u3_n172, 
       u2_u0_u3_n173, u2_u0_u3_n174, u2_u0_u3_n175, u2_u0_u3_n176, u2_u0_u3_n177, u2_u0_u3_n178, u2_u0_u3_n179, u2_u0_u3_n180, u2_u0_u3_n181, 
       u2_u0_u3_n182, u2_u0_u3_n183, u2_u0_u3_n184, u2_u0_u3_n185, u2_u0_u3_n186, u2_u0_u3_n94, u2_u0_u3_n95, u2_u0_u3_n96, u2_u0_u3_n97, 
       u2_u0_u3_n98, u2_u0_u3_n99, u2_u0_u4_n100, u2_u0_u4_n101, u2_u0_u4_n102, u2_u0_u4_n103, u2_u0_u4_n104, u2_u0_u4_n105, u2_u0_u4_n106, 
       u2_u0_u4_n107, u2_u0_u4_n108, u2_u0_u4_n109, u2_u0_u4_n110, u2_u0_u4_n111, u2_u0_u4_n112, u2_u0_u4_n113, u2_u0_u4_n114, u2_u0_u4_n115, 
       u2_u0_u4_n116, u2_u0_u4_n117, u2_u0_u4_n118, u2_u0_u4_n119, u2_u0_u4_n120, u2_u0_u4_n121, u2_u0_u4_n122, u2_u0_u4_n123, u2_u0_u4_n124, 
       u2_u0_u4_n125, u2_u0_u4_n126, u2_u0_u4_n127, u2_u0_u4_n128, u2_u0_u4_n129, u2_u0_u4_n130, u2_u0_u4_n131, u2_u0_u4_n132, u2_u0_u4_n133, 
       u2_u0_u4_n134, u2_u0_u4_n135, u2_u0_u4_n136, u2_u0_u4_n137, u2_u0_u4_n138, u2_u0_u4_n139, u2_u0_u4_n140, u2_u0_u4_n141, u2_u0_u4_n142, 
       u2_u0_u4_n143, u2_u0_u4_n144, u2_u0_u4_n145, u2_u0_u4_n146, u2_u0_u4_n147, u2_u0_u4_n148, u2_u0_u4_n149, u2_u0_u4_n150, u2_u0_u4_n151, 
       u2_u0_u4_n152, u2_u0_u4_n153, u2_u0_u4_n154, u2_u0_u4_n155, u2_u0_u4_n156, u2_u0_u4_n157, u2_u0_u4_n158, u2_u0_u4_n159, u2_u0_u4_n160, 
       u2_u0_u4_n161, u2_u0_u4_n162, u2_u0_u4_n163, u2_u0_u4_n164, u2_u0_u4_n165, u2_u0_u4_n166, u2_u0_u4_n167, u2_u0_u4_n168, u2_u0_u4_n169, 
       u2_u0_u4_n170, u2_u0_u4_n171, u2_u0_u4_n172, u2_u0_u4_n173, u2_u0_u4_n174, u2_u0_u4_n175, u2_u0_u4_n176, u2_u0_u4_n177, u2_u0_u4_n178, 
       u2_u0_u4_n179, u2_u0_u4_n180, u2_u0_u4_n181, u2_u0_u4_n182, u2_u0_u4_n183, u2_u0_u4_n184, u2_u0_u4_n185, u2_u0_u4_n186, u2_u0_u4_n94, 
       u2_u0_u4_n95, u2_u0_u4_n96, u2_u0_u4_n97, u2_u0_u4_n98, u2_u0_u4_n99, u2_u0_u5_n100, u2_u0_u5_n101, u2_u0_u5_n102, u2_u0_u5_n103, 
       u2_u0_u5_n104, u2_u0_u5_n105, u2_u0_u5_n106, u2_u0_u5_n107, u2_u0_u5_n108, u2_u0_u5_n109, u2_u0_u5_n110, u2_u0_u5_n111, u2_u0_u5_n112, 
       u2_u0_u5_n113, u2_u0_u5_n114, u2_u0_u5_n115, u2_u0_u5_n116, u2_u0_u5_n117, u2_u0_u5_n118, u2_u0_u5_n119, u2_u0_u5_n120, u2_u0_u5_n121, 
       u2_u0_u5_n122, u2_u0_u5_n123, u2_u0_u5_n124, u2_u0_u5_n125, u2_u0_u5_n126, u2_u0_u5_n127, u2_u0_u5_n128, u2_u0_u5_n129, u2_u0_u5_n130, 
       u2_u0_u5_n131, u2_u0_u5_n132, u2_u0_u5_n133, u2_u0_u5_n134, u2_u0_u5_n135, u2_u0_u5_n136, u2_u0_u5_n137, u2_u0_u5_n138, u2_u0_u5_n139, 
       u2_u0_u5_n140, u2_u0_u5_n141, u2_u0_u5_n142, u2_u0_u5_n143, u2_u0_u5_n144, u2_u0_u5_n145, u2_u0_u5_n146, u2_u0_u5_n147, u2_u0_u5_n148, 
       u2_u0_u5_n149, u2_u0_u5_n150, u2_u0_u5_n151, u2_u0_u5_n152, u2_u0_u5_n153, u2_u0_u5_n154, u2_u0_u5_n155, u2_u0_u5_n156, u2_u0_u5_n157, 
       u2_u0_u5_n158, u2_u0_u5_n159, u2_u0_u5_n160, u2_u0_u5_n161, u2_u0_u5_n162, u2_u0_u5_n163, u2_u0_u5_n164, u2_u0_u5_n165, u2_u0_u5_n166, 
       u2_u0_u5_n167, u2_u0_u5_n168, u2_u0_u5_n169, u2_u0_u5_n170, u2_u0_u5_n171, u2_u0_u5_n172, u2_u0_u5_n173, u2_u0_u5_n174, u2_u0_u5_n175, 
       u2_u0_u5_n176, u2_u0_u5_n177, u2_u0_u5_n178, u2_u0_u5_n179, u2_u0_u5_n180, u2_u0_u5_n181, u2_u0_u5_n182, u2_u0_u5_n183, u2_u0_u5_n184, 
       u2_u0_u5_n185, u2_u0_u5_n186, u2_u0_u5_n187, u2_u0_u5_n188, u2_u0_u5_n189, u2_u0_u5_n190, u2_u0_u5_n191, u2_u0_u5_n192, u2_u0_u5_n193, 
       u2_u0_u5_n194, u2_u0_u5_n195, u2_u0_u5_n196, u2_u0_u5_n99, u2_u0_u6_n100, u2_u0_u6_n101, u2_u0_u6_n102, u2_u0_u6_n103, u2_u0_u6_n104, 
       u2_u0_u6_n105, u2_u0_u6_n106, u2_u0_u6_n107, u2_u0_u6_n108, u2_u0_u6_n109, u2_u0_u6_n110, u2_u0_u6_n111, u2_u0_u6_n112, u2_u0_u6_n113, 
       u2_u0_u6_n114, u2_u0_u6_n115, u2_u0_u6_n116, u2_u0_u6_n117, u2_u0_u6_n118, u2_u0_u6_n119, u2_u0_u6_n120, u2_u0_u6_n121, u2_u0_u6_n122, 
       u2_u0_u6_n123, u2_u0_u6_n124, u2_u0_u6_n125, u2_u0_u6_n126, u2_u0_u6_n127, u2_u0_u6_n128, u2_u0_u6_n129, u2_u0_u6_n130, u2_u0_u6_n131, 
       u2_u0_u6_n132, u2_u0_u6_n133, u2_u0_u6_n134, u2_u0_u6_n135, u2_u0_u6_n136, u2_u0_u6_n137, u2_u0_u6_n138, u2_u0_u6_n139, u2_u0_u6_n140, 
       u2_u0_u6_n141, u2_u0_u6_n142, u2_u0_u6_n143, u2_u0_u6_n144, u2_u0_u6_n145, u2_u0_u6_n146, u2_u0_u6_n147, u2_u0_u6_n148, u2_u0_u6_n149, 
       u2_u0_u6_n150, u2_u0_u6_n151, u2_u0_u6_n152, u2_u0_u6_n153, u2_u0_u6_n154, u2_u0_u6_n155, u2_u0_u6_n156, u2_u0_u6_n157, u2_u0_u6_n158, 
       u2_u0_u6_n159, u2_u0_u6_n160, u2_u0_u6_n161, u2_u0_u6_n162, u2_u0_u6_n163, u2_u0_u6_n164, u2_u0_u6_n165, u2_u0_u6_n166, u2_u0_u6_n167, 
       u2_u0_u6_n168, u2_u0_u6_n169, u2_u0_u6_n170, u2_u0_u6_n171, u2_u0_u6_n172, u2_u0_u6_n173, u2_u0_u6_n174, u2_u0_u6_n88, u2_u0_u6_n89, 
       u2_u0_u6_n90, u2_u0_u6_n91, u2_u0_u6_n92, u2_u0_u6_n93, u2_u0_u6_n94, u2_u0_u6_n95, u2_u0_u6_n96, u2_u0_u6_n97, u2_u0_u6_n98, 
       u2_u0_u6_n99, u2_u0_u7_n100, u2_u0_u7_n101, u2_u0_u7_n102, u2_u0_u7_n103, u2_u0_u7_n104, u2_u0_u7_n105, u2_u0_u7_n106, u2_u0_u7_n107, 
       u2_u0_u7_n108, u2_u0_u7_n109, u2_u0_u7_n110, u2_u0_u7_n111, u2_u0_u7_n112, u2_u0_u7_n113, u2_u0_u7_n114, u2_u0_u7_n115, u2_u0_u7_n116, 
       u2_u0_u7_n117, u2_u0_u7_n118, u2_u0_u7_n119, u2_u0_u7_n120, u2_u0_u7_n121, u2_u0_u7_n122, u2_u0_u7_n123, u2_u0_u7_n124, u2_u0_u7_n125, 
       u2_u0_u7_n126, u2_u0_u7_n127, u2_u0_u7_n128, u2_u0_u7_n129, u2_u0_u7_n130, u2_u0_u7_n131, u2_u0_u7_n132, u2_u0_u7_n133, u2_u0_u7_n134, 
       u2_u0_u7_n135, u2_u0_u7_n136, u2_u0_u7_n137, u2_u0_u7_n138, u2_u0_u7_n139, u2_u0_u7_n140, u2_u0_u7_n141, u2_u0_u7_n142, u2_u0_u7_n143, 
       u2_u0_u7_n144, u2_u0_u7_n145, u2_u0_u7_n146, u2_u0_u7_n147, u2_u0_u7_n148, u2_u0_u7_n149, u2_u0_u7_n150, u2_u0_u7_n151, u2_u0_u7_n152, 
       u2_u0_u7_n153, u2_u0_u7_n154, u2_u0_u7_n155, u2_u0_u7_n156, u2_u0_u7_n157, u2_u0_u7_n158, u2_u0_u7_n159, u2_u0_u7_n160, u2_u0_u7_n161, 
       u2_u0_u7_n162, u2_u0_u7_n163, u2_u0_u7_n164, u2_u0_u7_n165, u2_u0_u7_n166, u2_u0_u7_n167, u2_u0_u7_n168, u2_u0_u7_n169, u2_u0_u7_n170, 
       u2_u0_u7_n171, u2_u0_u7_n172, u2_u0_u7_n173, u2_u0_u7_n174, u2_u0_u7_n175, u2_u0_u7_n176, u2_u0_u7_n177, u2_u0_u7_n178, u2_u0_u7_n179, 
       u2_u0_u7_n180, u2_u0_u7_n91, u2_u0_u7_n92, u2_u0_u7_n93, u2_u0_u7_n94, u2_u0_u7_n95, u2_u0_u7_n96, u2_u0_u7_n97, u2_u0_u7_n98, 
       u2_u0_u7_n99, u2_u11_X_1, u2_u11_X_10, u2_u11_X_11, u2_u11_X_12, u2_u11_X_2, u2_u11_X_3, u2_u11_X_4, u2_u11_X_5, 
       u2_u11_X_6, u2_u11_X_7, u2_u11_X_8, u2_u11_X_9, u2_u11_u0_n100, u2_u11_u0_n101, u2_u11_u0_n102, u2_u11_u0_n103, u2_u11_u0_n104, 
       u2_u11_u0_n105, u2_u11_u0_n106, u2_u11_u0_n107, u2_u11_u0_n108, u2_u11_u0_n109, u2_u11_u0_n110, u2_u11_u0_n111, u2_u11_u0_n112, u2_u11_u0_n113, 
       u2_u11_u0_n114, u2_u11_u0_n115, u2_u11_u0_n116, u2_u11_u0_n117, u2_u11_u0_n118, u2_u11_u0_n119, u2_u11_u0_n120, u2_u11_u0_n121, u2_u11_u0_n122, 
       u2_u11_u0_n123, u2_u11_u0_n124, u2_u11_u0_n125, u2_u11_u0_n126, u2_u11_u0_n127, u2_u11_u0_n128, u2_u11_u0_n129, u2_u11_u0_n130, u2_u11_u0_n131, 
       u2_u11_u0_n132, u2_u11_u0_n133, u2_u11_u0_n134, u2_u11_u0_n135, u2_u11_u0_n136, u2_u11_u0_n137, u2_u11_u0_n138, u2_u11_u0_n139, u2_u11_u0_n140, 
       u2_u11_u0_n141, u2_u11_u0_n142, u2_u11_u0_n143, u2_u11_u0_n144, u2_u11_u0_n145, u2_u11_u0_n146, u2_u11_u0_n147, u2_u11_u0_n148, u2_u11_u0_n149, 
       u2_u11_u0_n150, u2_u11_u0_n151, u2_u11_u0_n152, u2_u11_u0_n153, u2_u11_u0_n154, u2_u11_u0_n155, u2_u11_u0_n156, u2_u11_u0_n157, u2_u11_u0_n158, 
       u2_u11_u0_n159, u2_u11_u0_n160, u2_u11_u0_n161, u2_u11_u0_n162, u2_u11_u0_n163, u2_u11_u0_n164, u2_u11_u0_n165, u2_u11_u0_n166, u2_u11_u0_n167, 
       u2_u11_u0_n168, u2_u11_u0_n169, u2_u11_u0_n170, u2_u11_u0_n171, u2_u11_u0_n172, u2_u11_u0_n173, u2_u11_u0_n174, u2_u11_u0_n88, u2_u11_u0_n89, 
       u2_u11_u0_n90, u2_u11_u0_n91, u2_u11_u0_n92, u2_u11_u0_n93, u2_u11_u0_n94, u2_u11_u0_n95, u2_u11_u0_n96, u2_u11_u0_n97, u2_u11_u0_n98, 
       u2_u11_u0_n99, u2_u11_u1_n100, u2_u11_u1_n101, u2_u11_u1_n102, u2_u11_u1_n103, u2_u11_u1_n104, u2_u11_u1_n105, u2_u11_u1_n106, u2_u11_u1_n107, 
       u2_u11_u1_n108, u2_u11_u1_n109, u2_u11_u1_n110, u2_u11_u1_n111, u2_u11_u1_n112, u2_u11_u1_n113, u2_u11_u1_n114, u2_u11_u1_n115, u2_u11_u1_n116, 
       u2_u11_u1_n117, u2_u11_u1_n118, u2_u11_u1_n119, u2_u11_u1_n120, u2_u11_u1_n121, u2_u11_u1_n122, u2_u11_u1_n123, u2_u11_u1_n124, u2_u11_u1_n125, 
       u2_u11_u1_n126, u2_u11_u1_n127, u2_u11_u1_n128, u2_u11_u1_n129, u2_u11_u1_n130, u2_u11_u1_n131, u2_u11_u1_n132, u2_u11_u1_n133, u2_u11_u1_n134, 
       u2_u11_u1_n135, u2_u11_u1_n136, u2_u11_u1_n137, u2_u11_u1_n138, u2_u11_u1_n139, u2_u11_u1_n140, u2_u11_u1_n141, u2_u11_u1_n142, u2_u11_u1_n143, 
       u2_u11_u1_n144, u2_u11_u1_n145, u2_u11_u1_n146, u2_u11_u1_n147, u2_u11_u1_n148, u2_u11_u1_n149, u2_u11_u1_n150, u2_u11_u1_n151, u2_u11_u1_n152, 
       u2_u11_u1_n153, u2_u11_u1_n154, u2_u11_u1_n155, u2_u11_u1_n156, u2_u11_u1_n157, u2_u11_u1_n158, u2_u11_u1_n159, u2_u11_u1_n160, u2_u11_u1_n161, 
       u2_u11_u1_n162, u2_u11_u1_n163, u2_u11_u1_n164, u2_u11_u1_n165, u2_u11_u1_n166, u2_u11_u1_n167, u2_u11_u1_n168, u2_u11_u1_n169, u2_u11_u1_n170, 
       u2_u11_u1_n171, u2_u11_u1_n172, u2_u11_u1_n173, u2_u11_u1_n174, u2_u11_u1_n175, u2_u11_u1_n176, u2_u11_u1_n177, u2_u11_u1_n178, u2_u11_u1_n179, 
       u2_u11_u1_n180, u2_u11_u1_n181, u2_u11_u1_n182, u2_u11_u1_n183, u2_u11_u1_n184, u2_u11_u1_n185, u2_u11_u1_n186, u2_u11_u1_n187, u2_u11_u1_n188, 
       u2_u11_u1_n95, u2_u11_u1_n96, u2_u11_u1_n97, u2_u11_u1_n98, u2_u11_u1_n99, u2_u13_X_43, u2_u13_X_44, u2_u13_X_45, u2_u13_X_46, 
       u2_u13_X_47, u2_u13_X_48, u2_u13_u7_n100, u2_u13_u7_n101, u2_u13_u7_n102, u2_u13_u7_n103, u2_u13_u7_n104, u2_u13_u7_n105, u2_u13_u7_n106, 
       u2_u13_u7_n107, u2_u13_u7_n108, u2_u13_u7_n109, u2_u13_u7_n110, u2_u13_u7_n111, u2_u13_u7_n112, u2_u13_u7_n113, u2_u13_u7_n114, u2_u13_u7_n115, 
       u2_u13_u7_n116, u2_u13_u7_n117, u2_u13_u7_n118, u2_u13_u7_n119, u2_u13_u7_n120, u2_u13_u7_n121, u2_u13_u7_n122, u2_u13_u7_n123, u2_u13_u7_n124, 
       u2_u13_u7_n125, u2_u13_u7_n126, u2_u13_u7_n127, u2_u13_u7_n128, u2_u13_u7_n129, u2_u13_u7_n130, u2_u13_u7_n131, u2_u13_u7_n132, u2_u13_u7_n133, 
       u2_u13_u7_n134, u2_u13_u7_n135, u2_u13_u7_n136, u2_u13_u7_n137, u2_u13_u7_n138, u2_u13_u7_n139, u2_u13_u7_n140, u2_u13_u7_n141, u2_u13_u7_n142, 
       u2_u13_u7_n143, u2_u13_u7_n144, u2_u13_u7_n145, u2_u13_u7_n146, u2_u13_u7_n147, u2_u13_u7_n148, u2_u13_u7_n149, u2_u13_u7_n150, u2_u13_u7_n151, 
       u2_u13_u7_n152, u2_u13_u7_n153, u2_u13_u7_n154, u2_u13_u7_n155, u2_u13_u7_n156, u2_u13_u7_n157, u2_u13_u7_n158, u2_u13_u7_n159, u2_u13_u7_n160, 
       u2_u13_u7_n161, u2_u13_u7_n162, u2_u13_u7_n163, u2_u13_u7_n164, u2_u13_u7_n165, u2_u13_u7_n166, u2_u13_u7_n167, u2_u13_u7_n168, u2_u13_u7_n169, 
       u2_u13_u7_n170, u2_u13_u7_n171, u2_u13_u7_n172, u2_u13_u7_n173, u2_u13_u7_n174, u2_u13_u7_n175, u2_u13_u7_n176, u2_u13_u7_n177, u2_u13_u7_n178, 
       u2_u13_u7_n179, u2_u13_u7_n180, u2_u13_u7_n91, u2_u13_u7_n92, u2_u13_u7_n93, u2_u13_u7_n94, u2_u13_u7_n95, u2_u13_u7_n96, u2_u13_u7_n97, 
       u2_u13_u7_n98, u2_u13_u7_n99, u2_u1_X_31, u2_u1_X_32, u2_u1_X_33, u2_u1_X_34, u2_u1_X_35, u2_u1_X_36, u2_u1_X_37, 
       u2_u1_X_38, u2_u1_X_39, u2_u1_X_40, u2_u1_X_41, u2_u1_X_42, u2_u1_u5_n100, u2_u1_u5_n101, u2_u1_u5_n102, u2_u1_u5_n103, 
       u2_u1_u5_n104, u2_u1_u5_n105, u2_u1_u5_n106, u2_u1_u5_n107, u2_u1_u5_n108, u2_u1_u5_n109, u2_u1_u5_n110, u2_u1_u5_n111, u2_u1_u5_n112, 
       u2_u1_u5_n113, u2_u1_u5_n114, u2_u1_u5_n115, u2_u1_u5_n116, u2_u1_u5_n117, u2_u1_u5_n118, u2_u1_u5_n119, u2_u1_u5_n120, u2_u1_u5_n121, 
       u2_u1_u5_n122, u2_u1_u5_n123, u2_u1_u5_n124, u2_u1_u5_n125, u2_u1_u5_n126, u2_u1_u5_n127, u2_u1_u5_n128, u2_u1_u5_n129, u2_u1_u5_n130, 
       u2_u1_u5_n131, u2_u1_u5_n132, u2_u1_u5_n133, u2_u1_u5_n134, u2_u1_u5_n135, u2_u1_u5_n136, u2_u1_u5_n137, u2_u1_u5_n138, u2_u1_u5_n139, 
       u2_u1_u5_n140, u2_u1_u5_n141, u2_u1_u5_n142, u2_u1_u5_n143, u2_u1_u5_n144, u2_u1_u5_n145, u2_u1_u5_n146, u2_u1_u5_n147, u2_u1_u5_n148, 
       u2_u1_u5_n149, u2_u1_u5_n150, u2_u1_u5_n151, u2_u1_u5_n152, u2_u1_u5_n153, u2_u1_u5_n154, u2_u1_u5_n155, u2_u1_u5_n156, u2_u1_u5_n157, 
       u2_u1_u5_n158, u2_u1_u5_n159, u2_u1_u5_n160, u2_u1_u5_n161, u2_u1_u5_n162, u2_u1_u5_n163, u2_u1_u5_n164, u2_u1_u5_n165, u2_u1_u5_n166, 
       u2_u1_u5_n167, u2_u1_u5_n168, u2_u1_u5_n169, u2_u1_u5_n170, u2_u1_u5_n171, u2_u1_u5_n172, u2_u1_u5_n173, u2_u1_u5_n174, u2_u1_u5_n175, 
       u2_u1_u5_n176, u2_u1_u5_n177, u2_u1_u5_n178, u2_u1_u5_n179, u2_u1_u5_n180, u2_u1_u5_n181, u2_u1_u5_n182, u2_u1_u5_n183, u2_u1_u5_n184, 
       u2_u1_u5_n185, u2_u1_u5_n186, u2_u1_u5_n187, u2_u1_u5_n188, u2_u1_u5_n189, u2_u1_u5_n190, u2_u1_u5_n191, u2_u1_u5_n192, u2_u1_u5_n193, 
       u2_u1_u5_n194, u2_u1_u5_n195, u2_u1_u5_n196, u2_u1_u5_n99, u2_u1_u6_n100, u2_u1_u6_n101, u2_u1_u6_n102, u2_u1_u6_n103, u2_u1_u6_n104, 
       u2_u1_u6_n105, u2_u1_u6_n106, u2_u1_u6_n107, u2_u1_u6_n108, u2_u1_u6_n109, u2_u1_u6_n110, u2_u1_u6_n111, u2_u1_u6_n112, u2_u1_u6_n113, 
       u2_u1_u6_n114, u2_u1_u6_n115, u2_u1_u6_n116, u2_u1_u6_n117, u2_u1_u6_n118, u2_u1_u6_n119, u2_u1_u6_n120, u2_u1_u6_n121, u2_u1_u6_n122, 
       u2_u1_u6_n123, u2_u1_u6_n124, u2_u1_u6_n125, u2_u1_u6_n126, u2_u1_u6_n127, u2_u1_u6_n128, u2_u1_u6_n129, u2_u1_u6_n130, u2_u1_u6_n131, 
       u2_u1_u6_n132, u2_u1_u6_n133, u2_u1_u6_n134, u2_u1_u6_n135, u2_u1_u6_n136, u2_u1_u6_n137, u2_u1_u6_n138, u2_u1_u6_n139, u2_u1_u6_n140, 
       u2_u1_u6_n141, u2_u1_u6_n142, u2_u1_u6_n143, u2_u1_u6_n144, u2_u1_u6_n145, u2_u1_u6_n146, u2_u1_u6_n147, u2_u1_u6_n148, u2_u1_u6_n149, 
       u2_u1_u6_n150, u2_u1_u6_n151, u2_u1_u6_n152, u2_u1_u6_n153, u2_u1_u6_n154, u2_u1_u6_n155, u2_u1_u6_n156, u2_u1_u6_n157, u2_u1_u6_n158, 
       u2_u1_u6_n159, u2_u1_u6_n160, u2_u1_u6_n161, u2_u1_u6_n162, u2_u1_u6_n163, u2_u1_u6_n164, u2_u1_u6_n165, u2_u1_u6_n166, u2_u1_u6_n167, 
       u2_u1_u6_n168, u2_u1_u6_n169, u2_u1_u6_n170, u2_u1_u6_n171, u2_u1_u6_n172, u2_u1_u6_n173, u2_u1_u6_n174, u2_u1_u6_n88, u2_u1_u6_n89, 
       u2_u1_u6_n90, u2_u1_u6_n91, u2_u1_u6_n92, u2_u1_u6_n93, u2_u1_u6_n94, u2_u1_u6_n95, u2_u1_u6_n96, u2_u1_u6_n97, u2_u1_u6_n98, 
       u2_u1_u6_n99, u2_u4_X_1, u2_u4_X_10, u2_u4_X_11, u2_u4_X_12, u2_u4_X_13, u2_u4_X_14, u2_u4_X_15, u2_u4_X_16, 
       u2_u4_X_17, u2_u4_X_18, u2_u4_X_19, u2_u4_X_2, u2_u4_X_20, u2_u4_X_21, u2_u4_X_22, u2_u4_X_23, u2_u4_X_24, 
       u2_u4_X_25, u2_u4_X_26, u2_u4_X_27, u2_u4_X_28, u2_u4_X_29, u2_u4_X_3, u2_u4_X_30, u2_u4_X_4, u2_u4_X_5, 
       u2_u4_X_6, u2_u4_X_7, u2_u4_X_8, u2_u4_X_9, u2_u4_u0_n100, u2_u4_u0_n101, u2_u4_u0_n102, u2_u4_u0_n103, u2_u4_u0_n104, 
       u2_u4_u0_n105, u2_u4_u0_n106, u2_u4_u0_n107, u2_u4_u0_n108, u2_u4_u0_n109, u2_u4_u0_n110, u2_u4_u0_n111, u2_u4_u0_n112, u2_u4_u0_n113, 
       u2_u4_u0_n114, u2_u4_u0_n115, u2_u4_u0_n116, u2_u4_u0_n117, u2_u4_u0_n118, u2_u4_u0_n119, u2_u4_u0_n120, u2_u4_u0_n121, u2_u4_u0_n122, 
       u2_u4_u0_n123, u2_u4_u0_n124, u2_u4_u0_n125, u2_u4_u0_n126, u2_u4_u0_n127, u2_u4_u0_n128, u2_u4_u0_n129, u2_u4_u0_n130, u2_u4_u0_n131, 
       u2_u4_u0_n132, u2_u4_u0_n133, u2_u4_u0_n134, u2_u4_u0_n135, u2_u4_u0_n136, u2_u4_u0_n137, u2_u4_u0_n138, u2_u4_u0_n139, u2_u4_u0_n140, 
       u2_u4_u0_n141, u2_u4_u0_n142, u2_u4_u0_n143, u2_u4_u0_n144, u2_u4_u0_n145, u2_u4_u0_n146, u2_u4_u0_n147, u2_u4_u0_n148, u2_u4_u0_n149, 
       u2_u4_u0_n150, u2_u4_u0_n151, u2_u4_u0_n152, u2_u4_u0_n153, u2_u4_u0_n154, u2_u4_u0_n155, u2_u4_u0_n156, u2_u4_u0_n157, u2_u4_u0_n158, 
       u2_u4_u0_n159, u2_u4_u0_n160, u2_u4_u0_n161, u2_u4_u0_n162, u2_u4_u0_n163, u2_u4_u0_n164, u2_u4_u0_n165, u2_u4_u0_n166, u2_u4_u0_n167, 
       u2_u4_u0_n168, u2_u4_u0_n169, u2_u4_u0_n170, u2_u4_u0_n171, u2_u4_u0_n172, u2_u4_u0_n173, u2_u4_u0_n174, u2_u4_u0_n88, u2_u4_u0_n89, 
       u2_u4_u0_n90, u2_u4_u0_n91, u2_u4_u0_n92, u2_u4_u0_n93, u2_u4_u0_n94, u2_u4_u0_n95, u2_u4_u0_n96, u2_u4_u0_n97, u2_u4_u0_n98, 
       u2_u4_u0_n99, u2_u4_u1_n100, u2_u4_u1_n101, u2_u4_u1_n102, u2_u4_u1_n103, u2_u4_u1_n104, u2_u4_u1_n105, u2_u4_u1_n106, u2_u4_u1_n107, 
       u2_u4_u1_n108, u2_u4_u1_n109, u2_u4_u1_n110, u2_u4_u1_n111, u2_u4_u1_n112, u2_u4_u1_n113, u2_u4_u1_n114, u2_u4_u1_n115, u2_u4_u1_n116, 
       u2_u4_u1_n117, u2_u4_u1_n118, u2_u4_u1_n119, u2_u4_u1_n120, u2_u4_u1_n121, u2_u4_u1_n122, u2_u4_u1_n123, u2_u4_u1_n124, u2_u4_u1_n125, 
       u2_u4_u1_n126, u2_u4_u1_n127, u2_u4_u1_n128, u2_u4_u1_n129, u2_u4_u1_n130, u2_u4_u1_n131, u2_u4_u1_n132, u2_u4_u1_n133, u2_u4_u1_n134, 
       u2_u4_u1_n135, u2_u4_u1_n136, u2_u4_u1_n137, u2_u4_u1_n138, u2_u4_u1_n139, u2_u4_u1_n140, u2_u4_u1_n141, u2_u4_u1_n142, u2_u4_u1_n143, 
       u2_u4_u1_n144, u2_u4_u1_n145, u2_u4_u1_n146, u2_u4_u1_n147, u2_u4_u1_n148, u2_u4_u1_n149, u2_u4_u1_n150, u2_u4_u1_n151, u2_u4_u1_n152, 
       u2_u4_u1_n153, u2_u4_u1_n154, u2_u4_u1_n155, u2_u4_u1_n156, u2_u4_u1_n157, u2_u4_u1_n158, u2_u4_u1_n159, u2_u4_u1_n160, u2_u4_u1_n161, 
       u2_u4_u1_n162, u2_u4_u1_n163, u2_u4_u1_n164, u2_u4_u1_n165, u2_u4_u1_n166, u2_u4_u1_n167, u2_u4_u1_n168, u2_u4_u1_n169, u2_u4_u1_n170, 
       u2_u4_u1_n171, u2_u4_u1_n172, u2_u4_u1_n173, u2_u4_u1_n174, u2_u4_u1_n175, u2_u4_u1_n176, u2_u4_u1_n177, u2_u4_u1_n178, u2_u4_u1_n179, 
       u2_u4_u1_n180, u2_u4_u1_n181, u2_u4_u1_n182, u2_u4_u1_n183, u2_u4_u1_n184, u2_u4_u1_n185, u2_u4_u1_n186, u2_u4_u1_n187, u2_u4_u1_n188, 
       u2_u4_u1_n95, u2_u4_u1_n96, u2_u4_u1_n97, u2_u4_u1_n98, u2_u4_u1_n99, u2_u4_u2_n100, u2_u4_u2_n101, u2_u4_u2_n102, u2_u4_u2_n103, 
       u2_u4_u2_n104, u2_u4_u2_n105, u2_u4_u2_n106, u2_u4_u2_n107, u2_u4_u2_n108, u2_u4_u2_n109, u2_u4_u2_n110, u2_u4_u2_n111, u2_u4_u2_n112, 
       u2_u4_u2_n113, u2_u4_u2_n114, u2_u4_u2_n115, u2_u4_u2_n116, u2_u4_u2_n117, u2_u4_u2_n118, u2_u4_u2_n119, u2_u4_u2_n120, u2_u4_u2_n121, 
       u2_u4_u2_n122, u2_u4_u2_n123, u2_u4_u2_n124, u2_u4_u2_n125, u2_u4_u2_n126, u2_u4_u2_n127, u2_u4_u2_n128, u2_u4_u2_n129, u2_u4_u2_n130, 
       u2_u4_u2_n131, u2_u4_u2_n132, u2_u4_u2_n133, u2_u4_u2_n134, u2_u4_u2_n135, u2_u4_u2_n136, u2_u4_u2_n137, u2_u4_u2_n138, u2_u4_u2_n139, 
       u2_u4_u2_n140, u2_u4_u2_n141, u2_u4_u2_n142, u2_u4_u2_n143, u2_u4_u2_n144, u2_u4_u2_n145, u2_u4_u2_n146, u2_u4_u2_n147, u2_u4_u2_n148, 
       u2_u4_u2_n149, u2_u4_u2_n150, u2_u4_u2_n151, u2_u4_u2_n152, u2_u4_u2_n153, u2_u4_u2_n154, u2_u4_u2_n155, u2_u4_u2_n156, u2_u4_u2_n157, 
       u2_u4_u2_n158, u2_u4_u2_n159, u2_u4_u2_n160, u2_u4_u2_n161, u2_u4_u2_n162, u2_u4_u2_n163, u2_u4_u2_n164, u2_u4_u2_n165, u2_u4_u2_n166, 
       u2_u4_u2_n167, u2_u4_u2_n168, u2_u4_u2_n169, u2_u4_u2_n170, u2_u4_u2_n171, u2_u4_u2_n172, u2_u4_u2_n173, u2_u4_u2_n174, u2_u4_u2_n175, 
       u2_u4_u2_n176, u2_u4_u2_n177, u2_u4_u2_n178, u2_u4_u2_n179, u2_u4_u2_n180, u2_u4_u2_n181, u2_u4_u2_n182, u2_u4_u2_n183, u2_u4_u2_n184, 
       u2_u4_u2_n185, u2_u4_u2_n186, u2_u4_u2_n187, u2_u4_u2_n188, u2_u4_u2_n95, u2_u4_u2_n96, u2_u4_u2_n97, u2_u4_u2_n98, u2_u4_u2_n99, 
       u2_u4_u3_n100, u2_u4_u3_n101, u2_u4_u3_n102, u2_u4_u3_n103, u2_u4_u3_n104, u2_u4_u3_n105, u2_u4_u3_n106, u2_u4_u3_n107, u2_u4_u3_n108, 
       u2_u4_u3_n109, u2_u4_u3_n110, u2_u4_u3_n111, u2_u4_u3_n112, u2_u4_u3_n113, u2_u4_u3_n114, u2_u4_u3_n115, u2_u4_u3_n116, u2_u4_u3_n117, 
       u2_u4_u3_n118, u2_u4_u3_n119, u2_u4_u3_n120, u2_u4_u3_n121, u2_u4_u3_n122, u2_u4_u3_n123, u2_u4_u3_n124, u2_u4_u3_n125, u2_u4_u3_n126, 
       u2_u4_u3_n127, u2_u4_u3_n128, u2_u4_u3_n129, u2_u4_u3_n130, u2_u4_u3_n131, u2_u4_u3_n132, u2_u4_u3_n133, u2_u4_u3_n134, u2_u4_u3_n135, 
       u2_u4_u3_n136, u2_u4_u3_n137, u2_u4_u3_n138, u2_u4_u3_n139, u2_u4_u3_n140, u2_u4_u3_n141, u2_u4_u3_n142, u2_u4_u3_n143, u2_u4_u3_n144, 
       u2_u4_u3_n145, u2_u4_u3_n146, u2_u4_u3_n147, u2_u4_u3_n148, u2_u4_u3_n149, u2_u4_u3_n150, u2_u4_u3_n151, u2_u4_u3_n152, u2_u4_u3_n153, 
       u2_u4_u3_n154, u2_u4_u3_n155, u2_u4_u3_n156, u2_u4_u3_n157, u2_u4_u3_n158, u2_u4_u3_n159, u2_u4_u3_n160, u2_u4_u3_n161, u2_u4_u3_n162, 
       u2_u4_u3_n163, u2_u4_u3_n164, u2_u4_u3_n165, u2_u4_u3_n166, u2_u4_u3_n167, u2_u4_u3_n168, u2_u4_u3_n169, u2_u4_u3_n170, u2_u4_u3_n171, 
       u2_u4_u3_n172, u2_u4_u3_n173, u2_u4_u3_n174, u2_u4_u3_n175, u2_u4_u3_n176, u2_u4_u3_n177, u2_u4_u3_n178, u2_u4_u3_n179, u2_u4_u3_n180, 
       u2_u4_u3_n181, u2_u4_u3_n182, u2_u4_u3_n183, u2_u4_u3_n184, u2_u4_u3_n185, u2_u4_u3_n186, u2_u4_u3_n94, u2_u4_u3_n95, u2_u4_u3_n96, 
       u2_u4_u3_n97, u2_u4_u3_n98, u2_u4_u3_n99, u2_u4_u4_n100, u2_u4_u4_n101, u2_u4_u4_n102, u2_u4_u4_n103, u2_u4_u4_n104, u2_u4_u4_n105, 
       u2_u4_u4_n106, u2_u4_u4_n107, u2_u4_u4_n108, u2_u4_u4_n109, u2_u4_u4_n110, u2_u4_u4_n111, u2_u4_u4_n112, u2_u4_u4_n113, u2_u4_u4_n114, 
       u2_u4_u4_n115, u2_u4_u4_n116, u2_u4_u4_n117, u2_u4_u4_n118, u2_u4_u4_n119, u2_u4_u4_n120, u2_u4_u4_n121, u2_u4_u4_n122, u2_u4_u4_n123, 
       u2_u4_u4_n124, u2_u4_u4_n125, u2_u4_u4_n126, u2_u4_u4_n127, u2_u4_u4_n128, u2_u4_u4_n129, u2_u4_u4_n130, u2_u4_u4_n131, u2_u4_u4_n132, 
       u2_u4_u4_n133, u2_u4_u4_n134, u2_u4_u4_n135, u2_u4_u4_n136, u2_u4_u4_n137, u2_u4_u4_n138, u2_u4_u4_n139, u2_u4_u4_n140, u2_u4_u4_n141, 
       u2_u4_u4_n142, u2_u4_u4_n143, u2_u4_u4_n144, u2_u4_u4_n145, u2_u4_u4_n146, u2_u4_u4_n147, u2_u4_u4_n148, u2_u4_u4_n149, u2_u4_u4_n150, 
       u2_u4_u4_n151, u2_u4_u4_n152, u2_u4_u4_n153, u2_u4_u4_n154, u2_u4_u4_n155, u2_u4_u4_n156, u2_u4_u4_n157, u2_u4_u4_n158, u2_u4_u4_n159, 
       u2_u4_u4_n160, u2_u4_u4_n161, u2_u4_u4_n162, u2_u4_u4_n163, u2_u4_u4_n164, u2_u4_u4_n165, u2_u4_u4_n166, u2_u4_u4_n167, u2_u4_u4_n168, 
       u2_u4_u4_n169, u2_u4_u4_n170, u2_u4_u4_n171, u2_u4_u4_n172, u2_u4_u4_n173, u2_u4_u4_n174, u2_u4_u4_n175, u2_u4_u4_n176, u2_u4_u4_n177, 
       u2_u4_u4_n178, u2_u4_u4_n179, u2_u4_u4_n180, u2_u4_u4_n181, u2_u4_u4_n182, u2_u4_u4_n183, u2_u4_u4_n184, u2_u4_u4_n185, u2_u4_u4_n186, 
       u2_u4_u4_n94, u2_u4_u4_n95, u2_u4_u4_n96, u2_u4_u4_n97, u2_u4_u4_n98, u2_u4_u4_n99, u2_u7_X_1, u2_u7_X_13, u2_u7_X_14, 
       u2_u7_X_15, u2_u7_X_16, u2_u7_X_17, u2_u7_X_18, u2_u7_X_2, u2_u7_X_3, u2_u7_X_4, u2_u7_X_5, u2_u7_X_6, 
       u2_u7_u0_n100, u2_u7_u0_n101, u2_u7_u0_n102, u2_u7_u0_n103, u2_u7_u0_n104, u2_u7_u0_n105, u2_u7_u0_n106, u2_u7_u0_n107, u2_u7_u0_n108, 
       u2_u7_u0_n109, u2_u7_u0_n110, u2_u7_u0_n111, u2_u7_u0_n112, u2_u7_u0_n113, u2_u7_u0_n114, u2_u7_u0_n115, u2_u7_u0_n116, u2_u7_u0_n117, 
       u2_u7_u0_n118, u2_u7_u0_n119, u2_u7_u0_n120, u2_u7_u0_n121, u2_u7_u0_n122, u2_u7_u0_n123, u2_u7_u0_n124, u2_u7_u0_n125, u2_u7_u0_n126, 
       u2_u7_u0_n127, u2_u7_u0_n128, u2_u7_u0_n129, u2_u7_u0_n130, u2_u7_u0_n131, u2_u7_u0_n132, u2_u7_u0_n133, u2_u7_u0_n134, u2_u7_u0_n135, 
       u2_u7_u0_n136, u2_u7_u0_n137, u2_u7_u0_n138, u2_u7_u0_n139, u2_u7_u0_n140, u2_u7_u0_n141, u2_u7_u0_n142, u2_u7_u0_n143, u2_u7_u0_n144, 
       u2_u7_u0_n145, u2_u7_u0_n146, u2_u7_u0_n147, u2_u7_u0_n148, u2_u7_u0_n149, u2_u7_u0_n150, u2_u7_u0_n151, u2_u7_u0_n152, u2_u7_u0_n153, 
       u2_u7_u0_n154, u2_u7_u0_n155, u2_u7_u0_n156, u2_u7_u0_n157, u2_u7_u0_n158, u2_u7_u0_n159, u2_u7_u0_n160, u2_u7_u0_n161, u2_u7_u0_n162, 
       u2_u7_u0_n163, u2_u7_u0_n164, u2_u7_u0_n165, u2_u7_u0_n166, u2_u7_u0_n167, u2_u7_u0_n168, u2_u7_u0_n169, u2_u7_u0_n170, u2_u7_u0_n171, 
       u2_u7_u0_n172, u2_u7_u0_n173, u2_u7_u0_n174, u2_u7_u0_n88, u2_u7_u0_n89, u2_u7_u0_n90, u2_u7_u0_n91, u2_u7_u0_n92, u2_u7_u0_n93, 
       u2_u7_u0_n94, u2_u7_u0_n95, u2_u7_u0_n96, u2_u7_u0_n97, u2_u7_u0_n98, u2_u7_u0_n99, u2_u7_u2_n100, u2_u7_u2_n101, u2_u7_u2_n102, 
       u2_u7_u2_n103, u2_u7_u2_n104, u2_u7_u2_n105, u2_u7_u2_n106, u2_u7_u2_n107, u2_u7_u2_n108, u2_u7_u2_n109, u2_u7_u2_n110, u2_u7_u2_n111, 
       u2_u7_u2_n112, u2_u7_u2_n113, u2_u7_u2_n114, u2_u7_u2_n115, u2_u7_u2_n116, u2_u7_u2_n117, u2_u7_u2_n118, u2_u7_u2_n119, u2_u7_u2_n120, 
       u2_u7_u2_n121, u2_u7_u2_n122, u2_u7_u2_n123, u2_u7_u2_n124, u2_u7_u2_n125, u2_u7_u2_n126, u2_u7_u2_n127, u2_u7_u2_n128, u2_u7_u2_n129, 
       u2_u7_u2_n130, u2_u7_u2_n131, u2_u7_u2_n132, u2_u7_u2_n133, u2_u7_u2_n134, u2_u7_u2_n135, u2_u7_u2_n136, u2_u7_u2_n137, u2_u7_u2_n138, 
       u2_u7_u2_n139, u2_u7_u2_n140, u2_u7_u2_n141, u2_u7_u2_n142, u2_u7_u2_n143, u2_u7_u2_n144, u2_u7_u2_n145, u2_u7_u2_n146, u2_u7_u2_n147, 
       u2_u7_u2_n148, u2_u7_u2_n149, u2_u7_u2_n150, u2_u7_u2_n151, u2_u7_u2_n152, u2_u7_u2_n153, u2_u7_u2_n154, u2_u7_u2_n155, u2_u7_u2_n156, 
       u2_u7_u2_n157, u2_u7_u2_n158, u2_u7_u2_n159, u2_u7_u2_n160, u2_u7_u2_n161, u2_u7_u2_n162, u2_u7_u2_n163, u2_u7_u2_n164, u2_u7_u2_n165, 
       u2_u7_u2_n166, u2_u7_u2_n167, u2_u7_u2_n168, u2_u7_u2_n169, u2_u7_u2_n170, u2_u7_u2_n171, u2_u7_u2_n172, u2_u7_u2_n173, u2_u7_u2_n174, 
       u2_u7_u2_n175, u2_u7_u2_n176, u2_u7_u2_n177, u2_u7_u2_n178, u2_u7_u2_n179, u2_u7_u2_n180, u2_u7_u2_n181, u2_u7_u2_n182, u2_u7_u2_n183, 
       u2_u7_u2_n184, u2_u7_u2_n185, u2_u7_u2_n186, u2_u7_u2_n187, u2_u7_u2_n188, u2_u7_u2_n95, u2_u7_u2_n96, u2_u7_u2_n97, u2_u7_u2_n98, 
       u2_u7_u2_n99, u2_u8_X_19, u2_u8_X_20, u2_u8_X_21, u2_u8_X_22, u2_u8_X_23, u2_u8_X_24, u2_u8_X_25, u2_u8_X_26, 
       u2_u8_X_27, u2_u8_X_28, u2_u8_X_29, u2_u8_X_30, u2_u8_u3_n100, u2_u8_u3_n101, u2_u8_u3_n102, u2_u8_u3_n103, u2_u8_u3_n104, 
       u2_u8_u3_n105, u2_u8_u3_n106, u2_u8_u3_n107, u2_u8_u3_n108, u2_u8_u3_n109, u2_u8_u3_n110, u2_u8_u3_n111, u2_u8_u3_n112, u2_u8_u3_n113, 
       u2_u8_u3_n114, u2_u8_u3_n115, u2_u8_u3_n116, u2_u8_u3_n117, u2_u8_u3_n118, u2_u8_u3_n119, u2_u8_u3_n120, u2_u8_u3_n121, u2_u8_u3_n122, 
       u2_u8_u3_n123, u2_u8_u3_n124, u2_u8_u3_n125, u2_u8_u3_n126, u2_u8_u3_n127, u2_u8_u3_n128, u2_u8_u3_n129, u2_u8_u3_n130, u2_u8_u3_n131, 
       u2_u8_u3_n132, u2_u8_u3_n133, u2_u8_u3_n134, u2_u8_u3_n135, u2_u8_u3_n136, u2_u8_u3_n137, u2_u8_u3_n138, u2_u8_u3_n139, u2_u8_u3_n140, 
       u2_u8_u3_n141, u2_u8_u3_n142, u2_u8_u3_n143, u2_u8_u3_n144, u2_u8_u3_n145, u2_u8_u3_n146, u2_u8_u3_n147, u2_u8_u3_n148, u2_u8_u3_n149, 
       u2_u8_u3_n150, u2_u8_u3_n151, u2_u8_u3_n152, u2_u8_u3_n153, u2_u8_u3_n154, u2_u8_u3_n155, u2_u8_u3_n156, u2_u8_u3_n157, u2_u8_u3_n158, 
       u2_u8_u3_n159, u2_u8_u3_n160, u2_u8_u3_n161, u2_u8_u3_n162, u2_u8_u3_n163, u2_u8_u3_n164, u2_u8_u3_n165, u2_u8_u3_n166, u2_u8_u3_n167, 
       u2_u8_u3_n168, u2_u8_u3_n169, u2_u8_u3_n170, u2_u8_u3_n171, u2_u8_u3_n172, u2_u8_u3_n173, u2_u8_u3_n174, u2_u8_u3_n175, u2_u8_u3_n176, 
       u2_u8_u3_n177, u2_u8_u3_n178, u2_u8_u3_n179, u2_u8_u3_n180, u2_u8_u3_n181, u2_u8_u3_n182, u2_u8_u3_n183, u2_u8_u3_n184, u2_u8_u3_n185, 
       u2_u8_u3_n186, u2_u8_u3_n94, u2_u8_u3_n95, u2_u8_u3_n96, u2_u8_u3_n97, u2_u8_u3_n98, u2_u8_u3_n99, u2_u8_u4_n100, u2_u8_u4_n101, 
       u2_u8_u4_n102, u2_u8_u4_n103, u2_u8_u4_n104, u2_u8_u4_n105, u2_u8_u4_n106, u2_u8_u4_n107, u2_u8_u4_n108, u2_u8_u4_n109, u2_u8_u4_n110, 
       u2_u8_u4_n111, u2_u8_u4_n112, u2_u8_u4_n113, u2_u8_u4_n114, u2_u8_u4_n115, u2_u8_u4_n116, u2_u8_u4_n117, u2_u8_u4_n118, u2_u8_u4_n119, 
       u2_u8_u4_n120, u2_u8_u4_n121, u2_u8_u4_n122, u2_u8_u4_n123, u2_u8_u4_n124, u2_u8_u4_n125, u2_u8_u4_n126, u2_u8_u4_n127, u2_u8_u4_n128, 
       u2_u8_u4_n129, u2_u8_u4_n130, u2_u8_u4_n131, u2_u8_u4_n132, u2_u8_u4_n133, u2_u8_u4_n134, u2_u8_u4_n135, u2_u8_u4_n136, u2_u8_u4_n137, 
       u2_u8_u4_n138, u2_u8_u4_n139, u2_u8_u4_n140, u2_u8_u4_n141, u2_u8_u4_n142, u2_u8_u4_n143, u2_u8_u4_n144, u2_u8_u4_n145, u2_u8_u4_n146, 
       u2_u8_u4_n147, u2_u8_u4_n148, u2_u8_u4_n149, u2_u8_u4_n150, u2_u8_u4_n151, u2_u8_u4_n152, u2_u8_u4_n153, u2_u8_u4_n154, u2_u8_u4_n155, 
       u2_u8_u4_n156, u2_u8_u4_n157, u2_u8_u4_n158, u2_u8_u4_n159, u2_u8_u4_n160, u2_u8_u4_n161, u2_u8_u4_n162, u2_u8_u4_n163, u2_u8_u4_n164, 
       u2_u8_u4_n165, u2_u8_u4_n166, u2_u8_u4_n167, u2_u8_u4_n168, u2_u8_u4_n169, u2_u8_u4_n170, u2_u8_u4_n171, u2_u8_u4_n172, u2_u8_u4_n173, 
       u2_u8_u4_n174, u2_u8_u4_n175, u2_u8_u4_n176, u2_u8_u4_n177, u2_u8_u4_n178, u2_u8_u4_n179, u2_u8_u4_n180, u2_u8_u4_n181, u2_u8_u4_n182, 
       u2_u8_u4_n183, u2_u8_u4_n184, u2_u8_u4_n185, u2_u8_u4_n186, u2_u8_u4_n94, u2_u8_u4_n95, u2_u8_u4_n96, u2_u8_u4_n97, u2_u8_u4_n98, 
       u2_u8_u4_n99, u2_u9_X_31, u2_u9_X_32, u2_u9_X_33, u2_u9_X_34, u2_u9_X_35, u2_u9_X_36, u2_u9_X_37, u2_u9_X_38, 
       u2_u9_X_39, u2_u9_X_40, u2_u9_X_41, u2_u9_X_42, u2_u9_u5_n100, u2_u9_u5_n101, u2_u9_u5_n102, u2_u9_u5_n103, u2_u9_u5_n104, 
       u2_u9_u5_n105, u2_u9_u5_n106, u2_u9_u5_n107, u2_u9_u5_n108, u2_u9_u5_n109, u2_u9_u5_n110, u2_u9_u5_n111, u2_u9_u5_n112, u2_u9_u5_n113, 
       u2_u9_u5_n114, u2_u9_u5_n115, u2_u9_u5_n116, u2_u9_u5_n117, u2_u9_u5_n118, u2_u9_u5_n119, u2_u9_u5_n120, u2_u9_u5_n121, u2_u9_u5_n122, 
       u2_u9_u5_n123, u2_u9_u5_n124, u2_u9_u5_n125, u2_u9_u5_n126, u2_u9_u5_n127, u2_u9_u5_n128, u2_u9_u5_n129, u2_u9_u5_n130, u2_u9_u5_n131, 
       u2_u9_u5_n132, u2_u9_u5_n133, u2_u9_u5_n134, u2_u9_u5_n135, u2_u9_u5_n136, u2_u9_u5_n137, u2_u9_u5_n138, u2_u9_u5_n139, u2_u9_u5_n140, 
       u2_u9_u5_n141, u2_u9_u5_n142, u2_u9_u5_n143, u2_u9_u5_n144, u2_u9_u5_n145, u2_u9_u5_n146, u2_u9_u5_n147, u2_u9_u5_n148, u2_u9_u5_n149, 
       u2_u9_u5_n150, u2_u9_u5_n151, u2_u9_u5_n152, u2_u9_u5_n153, u2_u9_u5_n154, u2_u9_u5_n155, u2_u9_u5_n156, u2_u9_u5_n157, u2_u9_u5_n158, 
       u2_u9_u5_n159, u2_u9_u5_n160, u2_u9_u5_n161, u2_u9_u5_n162, u2_u9_u5_n163, u2_u9_u5_n164, u2_u9_u5_n165, u2_u9_u5_n166, u2_u9_u5_n167, 
       u2_u9_u5_n168, u2_u9_u5_n169, u2_u9_u5_n170, u2_u9_u5_n171, u2_u9_u5_n172, u2_u9_u5_n173, u2_u9_u5_n174, u2_u9_u5_n175, u2_u9_u5_n176, 
       u2_u9_u5_n177, u2_u9_u5_n178, u2_u9_u5_n179, u2_u9_u5_n180, u2_u9_u5_n181, u2_u9_u5_n182, u2_u9_u5_n183, u2_u9_u5_n184, u2_u9_u5_n185, 
       u2_u9_u5_n186, u2_u9_u5_n187, u2_u9_u5_n188, u2_u9_u5_n189, u2_u9_u5_n190, u2_u9_u5_n191, u2_u9_u5_n192, u2_u9_u5_n193, u2_u9_u5_n194, 
       u2_u9_u5_n195, u2_u9_u5_n196, u2_u9_u5_n99, u2_u9_u6_n100, u2_u9_u6_n101, u2_u9_u6_n102, u2_u9_u6_n103, u2_u9_u6_n104, u2_u9_u6_n105, 
       u2_u9_u6_n106, u2_u9_u6_n107, u2_u9_u6_n108, u2_u9_u6_n109, u2_u9_u6_n110, u2_u9_u6_n111, u2_u9_u6_n112, u2_u9_u6_n113, u2_u9_u6_n114, 
       u2_u9_u6_n115, u2_u9_u6_n116, u2_u9_u6_n117, u2_u9_u6_n118, u2_u9_u6_n119, u2_u9_u6_n120, u2_u9_u6_n121, u2_u9_u6_n122, u2_u9_u6_n123, 
       u2_u9_u6_n124, u2_u9_u6_n125, u2_u9_u6_n126, u2_u9_u6_n127, u2_u9_u6_n128, u2_u9_u6_n129, u2_u9_u6_n130, u2_u9_u6_n131, u2_u9_u6_n132, 
       u2_u9_u6_n133, u2_u9_u6_n134, u2_u9_u6_n135, u2_u9_u6_n136, u2_u9_u6_n137, u2_u9_u6_n138, u2_u9_u6_n139, u2_u9_u6_n140, u2_u9_u6_n141, 
       u2_u9_u6_n142, u2_u9_u6_n143, u2_u9_u6_n144, u2_u9_u6_n145, u2_u9_u6_n146, u2_u9_u6_n147, u2_u9_u6_n148, u2_u9_u6_n149, u2_u9_u6_n150, 
       u2_u9_u6_n151, u2_u9_u6_n152, u2_u9_u6_n153, u2_u9_u6_n154, u2_u9_u6_n155, u2_u9_u6_n156, u2_u9_u6_n157, u2_u9_u6_n158, u2_u9_u6_n159, 
       u2_u9_u6_n160, u2_u9_u6_n161, u2_u9_u6_n162, u2_u9_u6_n163, u2_u9_u6_n164, u2_u9_u6_n165, u2_u9_u6_n166, u2_u9_u6_n167, u2_u9_u6_n168, 
       u2_u9_u6_n169, u2_u9_u6_n170, u2_u9_u6_n171, u2_u9_u6_n172, u2_u9_u6_n173, u2_u9_u6_n174, u2_u9_u6_n88, u2_u9_u6_n89, u2_u9_u6_n90, 
       u2_u9_u6_n91, u2_u9_u6_n92, u2_u9_u6_n93, u2_u9_u6_n94, u2_u9_u6_n95, u2_u9_u6_n96, u2_u9_u6_n97, u2_u9_u6_n98, u2_u9_u6_n99, 
       u2_uk_n1000, u2_uk_n1041, u2_uk_n1055, u2_uk_n1057, u2_uk_n1099, u2_uk_n1101, u2_uk_n1110, u2_uk_n1124, u2_uk_n1126, 
       u2_uk_n1127, u2_uk_n1129, u2_uk_n1147, u2_uk_n1151, u2_uk_n1157, u2_uk_n1158, u2_uk_n1165, u2_uk_n1174, u2_uk_n291, 
       u2_uk_n294, u2_uk_n297, u2_uk_n301, u2_uk_n305, u2_uk_n306, u2_uk_n515, u2_uk_n518, u2_uk_n717, u2_uk_n930, 
       u2_uk_n973, u2_uk_n974, u2_uk_n975, u2_uk_n976, u2_uk_n977, u2_uk_n980, u2_uk_n981, u2_uk_n982, u2_uk_n985, 
       u2_uk_n987, u2_uk_n989,  u2_uk_n999;
  XOR2_X1 u0_U131 (.B( u0_L11_31 ) , .Z( u0_N414 ) , .A( u0_out12_31 ) );
  XOR2_X1 u0_U135 (.B( u0_L11_27 ) , .Z( u0_N410 ) , .A( u0_out12_27 ) );
  XOR2_X1 u0_U140 (.B( u0_L11_23 ) , .Z( u0_N406 ) , .A( u0_out12_23 ) );
  XOR2_X1 u0_U142 (.B( u0_L11_21 ) , .Z( u0_N404 ) , .A( u0_out12_21 ) );
  XOR2_X1 u0_U146 (.B( u0_L11_17 ) , .Z( u0_N400 ) , .A( u0_out12_17 ) );
  XOR2_X1 u0_U150 (.B( u0_L11_15 ) , .Z( u0_N398 ) , .A( u0_out12_15 ) );
  XOR2_X1 u0_U156 (.B( u0_L11_9 ) , .Z( u0_N392 ) , .A( u0_out12_9 ) );
  XOR2_X1 u0_U161 (.B( u0_L11_5 ) , .Z( u0_N388 ) , .A( u0_out12_5 ) );
  XOR2_X1 u0_U166 (.B( u0_L10_32 ) , .Z( u0_N383 ) , .A( u0_out11_32 ) );
  XOR2_X1 u0_U169 (.B( u0_L10_29 ) , .Z( u0_N380 ) , .A( u0_out11_29 ) );
  XOR2_X1 u0_U172 (.B( u0_L10_27 ) , .Z( u0_N378 ) , .A( u0_out11_27 ) );
  XOR2_X1 u0_U174 (.B( u0_L10_25 ) , .Z( u0_N376 ) , .A( u0_out11_25 ) );
  XOR2_X1 u0_U177 (.B( u0_L10_22 ) , .Z( u0_N373 ) , .A( u0_out11_22 ) );
  XOR2_X1 u0_U178 (.B( u0_L10_21 ) , .Z( u0_N372 ) , .A( u0_out11_21 ) );
  XOR2_X1 u0_U180 (.B( u0_L10_19 ) , .Z( u0_N370 ) , .A( u0_out11_19 ) );
  XOR2_X1 u0_U185 (.B( u0_L10_15 ) , .Z( u0_N366 ) , .A( u0_out11_15 ) );
  XOR2_X1 u0_U186 (.B( u0_L10_14 ) , .Z( u0_N365 ) , .A( u0_out11_14 ) );
  XOR2_X1 u0_U188 (.B( u0_L10_12 ) , .Z( u0_N363 ) , .A( u0_out11_12 ) );
  XOR2_X1 u0_U189 (.B( u0_L10_11 ) , .Z( u0_N362 ) , .A( u0_out11_11 ) );
  XOR2_X1 u0_U193 (.B( u0_L10_8 ) , .Z( u0_N359 ) , .A( u0_out11_8 ) );
  XOR2_X1 u0_U194 (.B( u0_L10_7 ) , .Z( u0_N358 ) , .A( u0_out11_7 ) );
  XOR2_X1 u0_U196 (.B( u0_L10_5 ) , .Z( u0_N356 ) , .A( u0_out11_5 ) );
  XOR2_X1 u0_U197 (.B( u0_L10_4 ) , .Z( u0_N355 ) , .A( u0_out11_4 ) );
  XOR2_X1 u0_U198 (.B( u0_L10_3 ) , .Z( u0_N354 ) , .A( u0_out11_3 ) );
  XOR2_X1 u0_U209 (.B( u0_L9_25 ) , .Z( u0_N344 ) , .A( u0_out10_25 ) );
  XOR2_X1 u0_U221 (.B( u0_L9_14 ) , .Z( u0_N333 ) , .A( u0_out10_14 ) );
  XOR2_X1 u0_U228 (.B( u0_L9_8 ) , .Z( u0_N327 ) , .A( u0_out10_8 ) );
  XOR2_X1 u0_U233 (.B( u0_L9_3 ) , .Z( u0_N322 ) , .A( u0_out10_3 ) );
  XOR2_X1 u0_u10_U26 (.B( u0_K11_30 ) , .A( u0_R9_21 ) , .Z( u0_u10_X_30 ) );
  XOR2_X1 u0_u10_U28 (.B( u0_K11_29 ) , .A( u0_R9_20 ) , .Z( u0_u10_X_29 ) );
  XOR2_X1 u0_u10_U29 (.B( u0_K11_28 ) , .A( u0_R9_19 ) , .Z( u0_u10_X_28 ) );
  XOR2_X1 u0_u10_U30 (.B( u0_K11_27 ) , .A( u0_R9_18 ) , .Z( u0_u10_X_27 ) );
  XOR2_X1 u0_u10_U31 (.B( u0_K11_26 ) , .A( u0_R9_17 ) , .Z( u0_u10_X_26 ) );
  XOR2_X1 u0_u10_U32 (.B( u0_K11_25 ) , .A( u0_R9_16 ) , .Z( u0_u10_X_25 ) );
  AOI21_X1 u0_u10_u4_U10 (.ZN( u0_u10_u4_n106 ) , .B2( u0_u10_u4_n146 ) , .B1( u0_u10_u4_n158 ) , .A( u0_u10_u4_n170 ) );
  AOI21_X1 u0_u10_u4_U11 (.ZN( u0_u10_u4_n108 ) , .B2( u0_u10_u4_n134 ) , .B1( u0_u10_u4_n155 ) , .A( u0_u10_u4_n156 ) );
  AOI21_X1 u0_u10_u4_U12 (.ZN( u0_u10_u4_n109 ) , .A( u0_u10_u4_n153 ) , .B1( u0_u10_u4_n159 ) , .B2( u0_u10_u4_n184 ) );
  AOI211_X1 u0_u10_u4_U13 (.B( u0_u10_u4_n136 ) , .A( u0_u10_u4_n137 ) , .C2( u0_u10_u4_n138 ) , .ZN( u0_u10_u4_n139 ) , .C1( u0_u10_u4_n182 ) );
  OAI22_X1 u0_u10_u4_U14 (.B2( u0_u10_u4_n135 ) , .ZN( u0_u10_u4_n137 ) , .B1( u0_u10_u4_n153 ) , .A1( u0_u10_u4_n155 ) , .A2( u0_u10_u4_n171 ) );
  AND3_X1 u0_u10_u4_U15 (.A2( u0_u10_u4_n134 ) , .ZN( u0_u10_u4_n135 ) , .A3( u0_u10_u4_n145 ) , .A1( u0_u10_u4_n157 ) );
  NAND2_X1 u0_u10_u4_U16 (.ZN( u0_u10_u4_n132 ) , .A2( u0_u10_u4_n170 ) , .A1( u0_u10_u4_n173 ) );
  AOI21_X1 u0_u10_u4_U17 (.B2( u0_u10_u4_n160 ) , .B1( u0_u10_u4_n161 ) , .ZN( u0_u10_u4_n162 ) , .A( u0_u10_u4_n170 ) );
  AOI21_X1 u0_u10_u4_U18 (.ZN( u0_u10_u4_n107 ) , .B2( u0_u10_u4_n143 ) , .A( u0_u10_u4_n174 ) , .B1( u0_u10_u4_n184 ) );
  AOI21_X1 u0_u10_u4_U19 (.B2( u0_u10_u4_n158 ) , .B1( u0_u10_u4_n159 ) , .ZN( u0_u10_u4_n163 ) , .A( u0_u10_u4_n174 ) );
  AOI21_X1 u0_u10_u4_U20 (.A( u0_u10_u4_n153 ) , .B2( u0_u10_u4_n154 ) , .B1( u0_u10_u4_n155 ) , .ZN( u0_u10_u4_n165 ) );
  AOI21_X1 u0_u10_u4_U21 (.A( u0_u10_u4_n156 ) , .B2( u0_u10_u4_n157 ) , .ZN( u0_u10_u4_n164 ) , .B1( u0_u10_u4_n184 ) );
  INV_X1 u0_u10_u4_U22 (.A( u0_u10_u4_n138 ) , .ZN( u0_u10_u4_n170 ) );
  AND2_X1 u0_u10_u4_U23 (.A2( u0_u10_u4_n120 ) , .ZN( u0_u10_u4_n155 ) , .A1( u0_u10_u4_n160 ) );
  INV_X1 u0_u10_u4_U24 (.A( u0_u10_u4_n156 ) , .ZN( u0_u10_u4_n175 ) );
  NAND2_X1 u0_u10_u4_U25 (.A2( u0_u10_u4_n118 ) , .ZN( u0_u10_u4_n131 ) , .A1( u0_u10_u4_n147 ) );
  NAND2_X1 u0_u10_u4_U26 (.A1( u0_u10_u4_n119 ) , .A2( u0_u10_u4_n120 ) , .ZN( u0_u10_u4_n130 ) );
  NAND2_X1 u0_u10_u4_U27 (.ZN( u0_u10_u4_n117 ) , .A2( u0_u10_u4_n118 ) , .A1( u0_u10_u4_n148 ) );
  NAND2_X1 u0_u10_u4_U28 (.ZN( u0_u10_u4_n129 ) , .A1( u0_u10_u4_n134 ) , .A2( u0_u10_u4_n148 ) );
  AND3_X1 u0_u10_u4_U29 (.A1( u0_u10_u4_n119 ) , .A2( u0_u10_u4_n143 ) , .A3( u0_u10_u4_n154 ) , .ZN( u0_u10_u4_n161 ) );
  NOR2_X1 u0_u10_u4_U3 (.ZN( u0_u10_u4_n121 ) , .A1( u0_u10_u4_n181 ) , .A2( u0_u10_u4_n182 ) );
  AND2_X1 u0_u10_u4_U30 (.A1( u0_u10_u4_n145 ) , .A2( u0_u10_u4_n147 ) , .ZN( u0_u10_u4_n159 ) );
  OR3_X1 u0_u10_u4_U31 (.A3( u0_u10_u4_n114 ) , .A2( u0_u10_u4_n115 ) , .A1( u0_u10_u4_n116 ) , .ZN( u0_u10_u4_n136 ) );
  AOI21_X1 u0_u10_u4_U32 (.A( u0_u10_u4_n113 ) , .ZN( u0_u10_u4_n116 ) , .B2( u0_u10_u4_n173 ) , .B1( u0_u10_u4_n174 ) );
  AOI21_X1 u0_u10_u4_U33 (.ZN( u0_u10_u4_n115 ) , .B2( u0_u10_u4_n145 ) , .B1( u0_u10_u4_n146 ) , .A( u0_u10_u4_n156 ) );
  OAI22_X1 u0_u10_u4_U34 (.ZN( u0_u10_u4_n114 ) , .A2( u0_u10_u4_n121 ) , .B1( u0_u10_u4_n160 ) , .B2( u0_u10_u4_n170 ) , .A1( u0_u10_u4_n171 ) );
  INV_X1 u0_u10_u4_U35 (.A( u0_u10_u4_n158 ) , .ZN( u0_u10_u4_n182 ) );
  INV_X1 u0_u10_u4_U36 (.ZN( u0_u10_u4_n181 ) , .A( u0_u10_u4_n96 ) );
  INV_X1 u0_u10_u4_U37 (.A( u0_u10_u4_n144 ) , .ZN( u0_u10_u4_n179 ) );
  INV_X1 u0_u10_u4_U38 (.A( u0_u10_u4_n157 ) , .ZN( u0_u10_u4_n178 ) );
  NAND2_X1 u0_u10_u4_U39 (.A2( u0_u10_u4_n154 ) , .A1( u0_u10_u4_n96 ) , .ZN( u0_u10_u4_n97 ) );
  INV_X1 u0_u10_u4_U4 (.A( u0_u10_u4_n117 ) , .ZN( u0_u10_u4_n184 ) );
  INV_X1 u0_u10_u4_U40 (.A( u0_u10_u4_n143 ) , .ZN( u0_u10_u4_n183 ) );
  NOR2_X1 u0_u10_u4_U41 (.ZN( u0_u10_u4_n138 ) , .A1( u0_u10_u4_n168 ) , .A2( u0_u10_u4_n169 ) );
  NOR2_X1 u0_u10_u4_U42 (.A1( u0_u10_u4_n150 ) , .A2( u0_u10_u4_n152 ) , .ZN( u0_u10_u4_n153 ) );
  NOR2_X1 u0_u10_u4_U43 (.A2( u0_u10_u4_n128 ) , .A1( u0_u10_u4_n138 ) , .ZN( u0_u10_u4_n156 ) );
  AOI22_X1 u0_u10_u4_U44 (.B2( u0_u10_u4_n122 ) , .A1( u0_u10_u4_n123 ) , .ZN( u0_u10_u4_n124 ) , .B1( u0_u10_u4_n128 ) , .A2( u0_u10_u4_n172 ) );
  INV_X1 u0_u10_u4_U45 (.A( u0_u10_u4_n153 ) , .ZN( u0_u10_u4_n172 ) );
  NAND2_X1 u0_u10_u4_U46 (.A2( u0_u10_u4_n120 ) , .ZN( u0_u10_u4_n123 ) , .A1( u0_u10_u4_n161 ) );
  AOI22_X1 u0_u10_u4_U47 (.B2( u0_u10_u4_n132 ) , .A2( u0_u10_u4_n133 ) , .ZN( u0_u10_u4_n140 ) , .A1( u0_u10_u4_n150 ) , .B1( u0_u10_u4_n179 ) );
  NAND2_X1 u0_u10_u4_U48 (.ZN( u0_u10_u4_n133 ) , .A2( u0_u10_u4_n146 ) , .A1( u0_u10_u4_n154 ) );
  NAND2_X1 u0_u10_u4_U49 (.A1( u0_u10_u4_n103 ) , .ZN( u0_u10_u4_n154 ) , .A2( u0_u10_u4_n98 ) );
  INV_X1 u0_u10_u4_U5 (.ZN( u0_u10_u4_n186 ) , .A( u0_u10_u4_n95 ) );
  NAND2_X1 u0_u10_u4_U50 (.A1( u0_u10_u4_n101 ) , .ZN( u0_u10_u4_n158 ) , .A2( u0_u10_u4_n99 ) );
  AOI21_X1 u0_u10_u4_U51 (.ZN( u0_u10_u4_n127 ) , .A( u0_u10_u4_n136 ) , .B2( u0_u10_u4_n150 ) , .B1( u0_u10_u4_n180 ) );
  INV_X1 u0_u10_u4_U52 (.A( u0_u10_u4_n160 ) , .ZN( u0_u10_u4_n180 ) );
  NAND2_X1 u0_u10_u4_U53 (.A2( u0_u10_u4_n104 ) , .A1( u0_u10_u4_n105 ) , .ZN( u0_u10_u4_n146 ) );
  NAND2_X1 u0_u10_u4_U54 (.A2( u0_u10_u4_n101 ) , .A1( u0_u10_u4_n102 ) , .ZN( u0_u10_u4_n160 ) );
  NAND2_X1 u0_u10_u4_U55 (.ZN( u0_u10_u4_n134 ) , .A1( u0_u10_u4_n98 ) , .A2( u0_u10_u4_n99 ) );
  NAND2_X1 u0_u10_u4_U56 (.A1( u0_u10_u4_n103 ) , .A2( u0_u10_u4_n104 ) , .ZN( u0_u10_u4_n143 ) );
  NAND2_X1 u0_u10_u4_U57 (.A2( u0_u10_u4_n105 ) , .ZN( u0_u10_u4_n145 ) , .A1( u0_u10_u4_n98 ) );
  NAND2_X1 u0_u10_u4_U58 (.A1( u0_u10_u4_n100 ) , .A2( u0_u10_u4_n105 ) , .ZN( u0_u10_u4_n120 ) );
  NAND2_X1 u0_u10_u4_U59 (.A1( u0_u10_u4_n102 ) , .A2( u0_u10_u4_n104 ) , .ZN( u0_u10_u4_n148 ) );
  OAI221_X1 u0_u10_u4_U6 (.C1( u0_u10_u4_n134 ) , .B1( u0_u10_u4_n158 ) , .B2( u0_u10_u4_n171 ) , .C2( u0_u10_u4_n173 ) , .A( u0_u10_u4_n94 ) , .ZN( u0_u10_u4_n95 ) );
  NAND2_X1 u0_u10_u4_U60 (.A2( u0_u10_u4_n100 ) , .A1( u0_u10_u4_n103 ) , .ZN( u0_u10_u4_n157 ) );
  INV_X1 u0_u10_u4_U61 (.A( u0_u10_u4_n150 ) , .ZN( u0_u10_u4_n173 ) );
  INV_X1 u0_u10_u4_U62 (.A( u0_u10_u4_n152 ) , .ZN( u0_u10_u4_n171 ) );
  NAND2_X1 u0_u10_u4_U63 (.A1( u0_u10_u4_n100 ) , .ZN( u0_u10_u4_n118 ) , .A2( u0_u10_u4_n99 ) );
  NAND2_X1 u0_u10_u4_U64 (.A2( u0_u10_u4_n100 ) , .A1( u0_u10_u4_n102 ) , .ZN( u0_u10_u4_n144 ) );
  NAND2_X1 u0_u10_u4_U65 (.A2( u0_u10_u4_n101 ) , .A1( u0_u10_u4_n105 ) , .ZN( u0_u10_u4_n96 ) );
  INV_X1 u0_u10_u4_U66 (.A( u0_u10_u4_n128 ) , .ZN( u0_u10_u4_n174 ) );
  NAND2_X1 u0_u10_u4_U67 (.A2( u0_u10_u4_n102 ) , .ZN( u0_u10_u4_n119 ) , .A1( u0_u10_u4_n98 ) );
  NAND2_X1 u0_u10_u4_U68 (.A2( u0_u10_u4_n101 ) , .A1( u0_u10_u4_n103 ) , .ZN( u0_u10_u4_n147 ) );
  NAND2_X1 u0_u10_u4_U69 (.A2( u0_u10_u4_n104 ) , .ZN( u0_u10_u4_n113 ) , .A1( u0_u10_u4_n99 ) );
  AOI222_X1 u0_u10_u4_U7 (.B2( u0_u10_u4_n132 ) , .A1( u0_u10_u4_n138 ) , .C2( u0_u10_u4_n175 ) , .A2( u0_u10_u4_n179 ) , .C1( u0_u10_u4_n181 ) , .B1( u0_u10_u4_n185 ) , .ZN( u0_u10_u4_n94 ) );
  NOR2_X1 u0_u10_u4_U70 (.A2( u0_u10_X_28 ) , .ZN( u0_u10_u4_n150 ) , .A1( u0_u10_u4_n168 ) );
  NOR2_X1 u0_u10_u4_U71 (.A2( u0_u10_X_29 ) , .ZN( u0_u10_u4_n152 ) , .A1( u0_u10_u4_n169 ) );
  NOR2_X1 u0_u10_u4_U72 (.A2( u0_u10_X_30 ) , .ZN( u0_u10_u4_n105 ) , .A1( u0_u10_u4_n176 ) );
  NOR2_X1 u0_u10_u4_U73 (.A2( u0_u10_X_26 ) , .ZN( u0_u10_u4_n100 ) , .A1( u0_u10_u4_n177 ) );
  NOR2_X1 u0_u10_u4_U74 (.A2( u0_u10_X_28 ) , .A1( u0_u10_X_29 ) , .ZN( u0_u10_u4_n128 ) );
  NOR2_X1 u0_u10_u4_U75 (.A2( u0_u10_X_27 ) , .A1( u0_u10_X_30 ) , .ZN( u0_u10_u4_n102 ) );
  NOR2_X1 u0_u10_u4_U76 (.A2( u0_u10_X_25 ) , .A1( u0_u10_X_26 ) , .ZN( u0_u10_u4_n98 ) );
  AND2_X1 u0_u10_u4_U77 (.A2( u0_u10_X_25 ) , .A1( u0_u10_X_26 ) , .ZN( u0_u10_u4_n104 ) );
  AND2_X1 u0_u10_u4_U78 (.A1( u0_u10_X_30 ) , .A2( u0_u10_u4_n176 ) , .ZN( u0_u10_u4_n99 ) );
  AND2_X1 u0_u10_u4_U79 (.A1( u0_u10_X_26 ) , .ZN( u0_u10_u4_n101 ) , .A2( u0_u10_u4_n177 ) );
  INV_X1 u0_u10_u4_U8 (.A( u0_u10_u4_n113 ) , .ZN( u0_u10_u4_n185 ) );
  AND2_X1 u0_u10_u4_U80 (.A1( u0_u10_X_27 ) , .A2( u0_u10_X_30 ) , .ZN( u0_u10_u4_n103 ) );
  INV_X1 u0_u10_u4_U81 (.A( u0_u10_X_28 ) , .ZN( u0_u10_u4_n169 ) );
  INV_X1 u0_u10_u4_U82 (.A( u0_u10_X_29 ) , .ZN( u0_u10_u4_n168 ) );
  INV_X1 u0_u10_u4_U83 (.A( u0_u10_X_25 ) , .ZN( u0_u10_u4_n177 ) );
  INV_X1 u0_u10_u4_U84 (.A( u0_u10_X_27 ) , .ZN( u0_u10_u4_n176 ) );
  NAND4_X1 u0_u10_u4_U85 (.ZN( u0_out10_25 ) , .A4( u0_u10_u4_n139 ) , .A3( u0_u10_u4_n140 ) , .A2( u0_u10_u4_n141 ) , .A1( u0_u10_u4_n142 ) );
  OAI21_X1 u0_u10_u4_U86 (.A( u0_u10_u4_n128 ) , .B2( u0_u10_u4_n129 ) , .B1( u0_u10_u4_n130 ) , .ZN( u0_u10_u4_n142 ) );
  OAI21_X1 u0_u10_u4_U87 (.B2( u0_u10_u4_n131 ) , .ZN( u0_u10_u4_n141 ) , .A( u0_u10_u4_n175 ) , .B1( u0_u10_u4_n183 ) );
  NAND4_X1 u0_u10_u4_U88 (.ZN( u0_out10_14 ) , .A4( u0_u10_u4_n124 ) , .A3( u0_u10_u4_n125 ) , .A2( u0_u10_u4_n126 ) , .A1( u0_u10_u4_n127 ) );
  AOI22_X1 u0_u10_u4_U89 (.B2( u0_u10_u4_n117 ) , .ZN( u0_u10_u4_n126 ) , .A1( u0_u10_u4_n129 ) , .B1( u0_u10_u4_n152 ) , .A2( u0_u10_u4_n175 ) );
  NOR4_X1 u0_u10_u4_U9 (.A4( u0_u10_u4_n106 ) , .A3( u0_u10_u4_n107 ) , .A2( u0_u10_u4_n108 ) , .A1( u0_u10_u4_n109 ) , .ZN( u0_u10_u4_n110 ) );
  AOI22_X1 u0_u10_u4_U90 (.ZN( u0_u10_u4_n125 ) , .B2( u0_u10_u4_n131 ) , .A2( u0_u10_u4_n132 ) , .B1( u0_u10_u4_n138 ) , .A1( u0_u10_u4_n178 ) );
  NAND4_X1 u0_u10_u4_U91 (.ZN( u0_out10_8 ) , .A4( u0_u10_u4_n110 ) , .A3( u0_u10_u4_n111 ) , .A2( u0_u10_u4_n112 ) , .A1( u0_u10_u4_n186 ) );
  NAND2_X1 u0_u10_u4_U92 (.ZN( u0_u10_u4_n112 ) , .A2( u0_u10_u4_n130 ) , .A1( u0_u10_u4_n150 ) );
  AOI22_X1 u0_u10_u4_U93 (.ZN( u0_u10_u4_n111 ) , .B2( u0_u10_u4_n132 ) , .A1( u0_u10_u4_n152 ) , .B1( u0_u10_u4_n178 ) , .A2( u0_u10_u4_n97 ) );
  AOI22_X1 u0_u10_u4_U94 (.B2( u0_u10_u4_n149 ) , .B1( u0_u10_u4_n150 ) , .A2( u0_u10_u4_n151 ) , .A1( u0_u10_u4_n152 ) , .ZN( u0_u10_u4_n167 ) );
  NOR4_X1 u0_u10_u4_U95 (.A4( u0_u10_u4_n162 ) , .A3( u0_u10_u4_n163 ) , .A2( u0_u10_u4_n164 ) , .A1( u0_u10_u4_n165 ) , .ZN( u0_u10_u4_n166 ) );
  NAND3_X1 u0_u10_u4_U96 (.ZN( u0_out10_3 ) , .A3( u0_u10_u4_n166 ) , .A1( u0_u10_u4_n167 ) , .A2( u0_u10_u4_n186 ) );
  NAND3_X1 u0_u10_u4_U97 (.A3( u0_u10_u4_n146 ) , .A2( u0_u10_u4_n147 ) , .A1( u0_u10_u4_n148 ) , .ZN( u0_u10_u4_n149 ) );
  NAND3_X1 u0_u10_u4_U98 (.A3( u0_u10_u4_n143 ) , .A2( u0_u10_u4_n144 ) , .A1( u0_u10_u4_n145 ) , .ZN( u0_u10_u4_n151 ) );
  NAND3_X1 u0_u10_u4_U99 (.A3( u0_u10_u4_n121 ) , .ZN( u0_u10_u4_n122 ) , .A2( u0_u10_u4_n144 ) , .A1( u0_u10_u4_n154 ) );
  XOR2_X1 u0_u11_U10 (.B( u0_K12_45 ) , .A( u0_R10_30 ) , .Z( u0_u11_X_45 ) );
  XOR2_X1 u0_u11_U11 (.B( u0_K12_44 ) , .A( u0_R10_29 ) , .Z( u0_u11_X_44 ) );
  XOR2_X1 u0_u11_U12 (.B( u0_K12_43 ) , .A( u0_R10_28 ) , .Z( u0_u11_X_43 ) );
  XOR2_X1 u0_u11_U13 (.B( u0_K12_42 ) , .A( u0_R10_29 ) , .Z( u0_u11_X_42 ) );
  XOR2_X1 u0_u11_U14 (.B( u0_K12_41 ) , .A( u0_R10_28 ) , .Z( u0_u11_X_41 ) );
  XOR2_X1 u0_u11_U15 (.B( u0_K12_40 ) , .A( u0_R10_27 ) , .Z( u0_u11_X_40 ) );
  XOR2_X1 u0_u11_U17 (.B( u0_K12_39 ) , .A( u0_R10_26 ) , .Z( u0_u11_X_39 ) );
  XOR2_X1 u0_u11_U18 (.B( u0_K12_38 ) , .A( u0_R10_25 ) , .Z( u0_u11_X_38 ) );
  XOR2_X1 u0_u11_U19 (.B( u0_K12_37 ) , .A( u0_R10_24 ) , .Z( u0_u11_X_37 ) );
  XOR2_X1 u0_u11_U20 (.B( u0_K12_36 ) , .A( u0_R10_25 ) , .Z( u0_u11_X_36 ) );
  XOR2_X1 u0_u11_U21 (.B( u0_K12_35 ) , .A( u0_R10_24 ) , .Z( u0_u11_X_35 ) );
  XOR2_X1 u0_u11_U22 (.B( u0_K12_34 ) , .A( u0_R10_23 ) , .Z( u0_u11_X_34 ) );
  XOR2_X1 u0_u11_U23 (.B( u0_K12_33 ) , .A( u0_R10_22 ) , .Z( u0_u11_X_33 ) );
  XOR2_X1 u0_u11_U24 (.B( u0_K12_32 ) , .A( u0_R10_21 ) , .Z( u0_u11_X_32 ) );
  XOR2_X1 u0_u11_U25 (.B( u0_K12_31 ) , .A( u0_R10_20 ) , .Z( u0_u11_X_31 ) );
  XOR2_X1 u0_u11_U26 (.B( u0_K12_30 ) , .A( u0_R10_21 ) , .Z( u0_u11_X_30 ) );
  XOR2_X1 u0_u11_U28 (.B( u0_K12_29 ) , .A( u0_R10_20 ) , .Z( u0_u11_X_29 ) );
  XOR2_X1 u0_u11_U29 (.B( u0_K12_28 ) , .A( u0_R10_19 ) , .Z( u0_u11_X_28 ) );
  XOR2_X1 u0_u11_U30 (.B( u0_K12_27 ) , .A( u0_R10_18 ) , .Z( u0_u11_X_27 ) );
  XOR2_X1 u0_u11_U31 (.B( u0_K12_26 ) , .A( u0_R10_17 ) , .Z( u0_u11_X_26 ) );
  XOR2_X1 u0_u11_U32 (.B( u0_K12_25 ) , .A( u0_R10_16 ) , .Z( u0_u11_X_25 ) );
  XOR2_X1 u0_u11_U7 (.B( u0_K12_48 ) , .A( u0_R10_1 ) , .Z( u0_u11_X_48 ) );
  XOR2_X1 u0_u11_U8 (.B( u0_K12_47 ) , .A( u0_R10_32 ) , .Z( u0_u11_X_47 ) );
  XOR2_X1 u0_u11_U9 (.B( u0_K12_46 ) , .A( u0_R10_31 ) , .Z( u0_u11_X_46 ) );
  OAI22_X1 u0_u11_u4_U10 (.B2( u0_u11_u4_n135 ) , .ZN( u0_u11_u4_n137 ) , .B1( u0_u11_u4_n153 ) , .A1( u0_u11_u4_n155 ) , .A2( u0_u11_u4_n171 ) );
  AND3_X1 u0_u11_u4_U11 (.A2( u0_u11_u4_n134 ) , .ZN( u0_u11_u4_n135 ) , .A3( u0_u11_u4_n145 ) , .A1( u0_u11_u4_n157 ) );
  NAND2_X1 u0_u11_u4_U12 (.ZN( u0_u11_u4_n132 ) , .A2( u0_u11_u4_n170 ) , .A1( u0_u11_u4_n173 ) );
  AOI21_X1 u0_u11_u4_U13 (.B2( u0_u11_u4_n160 ) , .B1( u0_u11_u4_n161 ) , .ZN( u0_u11_u4_n162 ) , .A( u0_u11_u4_n170 ) );
  AOI21_X1 u0_u11_u4_U14 (.ZN( u0_u11_u4_n107 ) , .B2( u0_u11_u4_n143 ) , .A( u0_u11_u4_n174 ) , .B1( u0_u11_u4_n184 ) );
  AOI21_X1 u0_u11_u4_U15 (.B2( u0_u11_u4_n158 ) , .B1( u0_u11_u4_n159 ) , .ZN( u0_u11_u4_n163 ) , .A( u0_u11_u4_n174 ) );
  AOI21_X1 u0_u11_u4_U16 (.A( u0_u11_u4_n153 ) , .B2( u0_u11_u4_n154 ) , .B1( u0_u11_u4_n155 ) , .ZN( u0_u11_u4_n165 ) );
  AOI21_X1 u0_u11_u4_U17 (.A( u0_u11_u4_n156 ) , .B2( u0_u11_u4_n157 ) , .ZN( u0_u11_u4_n164 ) , .B1( u0_u11_u4_n184 ) );
  INV_X1 u0_u11_u4_U18 (.A( u0_u11_u4_n138 ) , .ZN( u0_u11_u4_n170 ) );
  AND2_X1 u0_u11_u4_U19 (.A2( u0_u11_u4_n120 ) , .ZN( u0_u11_u4_n155 ) , .A1( u0_u11_u4_n160 ) );
  INV_X1 u0_u11_u4_U20 (.A( u0_u11_u4_n156 ) , .ZN( u0_u11_u4_n175 ) );
  NAND2_X1 u0_u11_u4_U21 (.A2( u0_u11_u4_n118 ) , .ZN( u0_u11_u4_n131 ) , .A1( u0_u11_u4_n147 ) );
  NAND2_X1 u0_u11_u4_U22 (.A1( u0_u11_u4_n119 ) , .A2( u0_u11_u4_n120 ) , .ZN( u0_u11_u4_n130 ) );
  NAND2_X1 u0_u11_u4_U23 (.ZN( u0_u11_u4_n117 ) , .A2( u0_u11_u4_n118 ) , .A1( u0_u11_u4_n148 ) );
  NAND2_X1 u0_u11_u4_U24 (.ZN( u0_u11_u4_n129 ) , .A1( u0_u11_u4_n134 ) , .A2( u0_u11_u4_n148 ) );
  AND3_X1 u0_u11_u4_U25 (.A1( u0_u11_u4_n119 ) , .A2( u0_u11_u4_n143 ) , .A3( u0_u11_u4_n154 ) , .ZN( u0_u11_u4_n161 ) );
  AND2_X1 u0_u11_u4_U26 (.A1( u0_u11_u4_n145 ) , .A2( u0_u11_u4_n147 ) , .ZN( u0_u11_u4_n159 ) );
  OR3_X1 u0_u11_u4_U27 (.A3( u0_u11_u4_n114 ) , .A2( u0_u11_u4_n115 ) , .A1( u0_u11_u4_n116 ) , .ZN( u0_u11_u4_n136 ) );
  AOI21_X1 u0_u11_u4_U28 (.A( u0_u11_u4_n113 ) , .ZN( u0_u11_u4_n116 ) , .B2( u0_u11_u4_n173 ) , .B1( u0_u11_u4_n174 ) );
  AOI21_X1 u0_u11_u4_U29 (.ZN( u0_u11_u4_n115 ) , .B2( u0_u11_u4_n145 ) , .B1( u0_u11_u4_n146 ) , .A( u0_u11_u4_n156 ) );
  NOR2_X1 u0_u11_u4_U3 (.ZN( u0_u11_u4_n121 ) , .A1( u0_u11_u4_n181 ) , .A2( u0_u11_u4_n182 ) );
  OAI22_X1 u0_u11_u4_U30 (.ZN( u0_u11_u4_n114 ) , .A2( u0_u11_u4_n121 ) , .B1( u0_u11_u4_n160 ) , .B2( u0_u11_u4_n170 ) , .A1( u0_u11_u4_n171 ) );
  INV_X1 u0_u11_u4_U31 (.A( u0_u11_u4_n158 ) , .ZN( u0_u11_u4_n182 ) );
  INV_X1 u0_u11_u4_U32 (.ZN( u0_u11_u4_n181 ) , .A( u0_u11_u4_n96 ) );
  INV_X1 u0_u11_u4_U33 (.A( u0_u11_u4_n144 ) , .ZN( u0_u11_u4_n179 ) );
  INV_X1 u0_u11_u4_U34 (.A( u0_u11_u4_n157 ) , .ZN( u0_u11_u4_n178 ) );
  NAND2_X1 u0_u11_u4_U35 (.A2( u0_u11_u4_n154 ) , .A1( u0_u11_u4_n96 ) , .ZN( u0_u11_u4_n97 ) );
  INV_X1 u0_u11_u4_U36 (.ZN( u0_u11_u4_n186 ) , .A( u0_u11_u4_n95 ) );
  OAI221_X1 u0_u11_u4_U37 (.C1( u0_u11_u4_n134 ) , .B1( u0_u11_u4_n158 ) , .B2( u0_u11_u4_n171 ) , .C2( u0_u11_u4_n173 ) , .A( u0_u11_u4_n94 ) , .ZN( u0_u11_u4_n95 ) );
  AOI222_X1 u0_u11_u4_U38 (.B2( u0_u11_u4_n132 ) , .A1( u0_u11_u4_n138 ) , .C2( u0_u11_u4_n175 ) , .A2( u0_u11_u4_n179 ) , .C1( u0_u11_u4_n181 ) , .B1( u0_u11_u4_n185 ) , .ZN( u0_u11_u4_n94 ) );
  INV_X1 u0_u11_u4_U39 (.A( u0_u11_u4_n113 ) , .ZN( u0_u11_u4_n185 ) );
  INV_X1 u0_u11_u4_U4 (.A( u0_u11_u4_n117 ) , .ZN( u0_u11_u4_n184 ) );
  INV_X1 u0_u11_u4_U40 (.A( u0_u11_u4_n143 ) , .ZN( u0_u11_u4_n183 ) );
  NOR2_X1 u0_u11_u4_U41 (.ZN( u0_u11_u4_n138 ) , .A1( u0_u11_u4_n168 ) , .A2( u0_u11_u4_n169 ) );
  NOR2_X1 u0_u11_u4_U42 (.A1( u0_u11_u4_n150 ) , .A2( u0_u11_u4_n152 ) , .ZN( u0_u11_u4_n153 ) );
  NOR2_X1 u0_u11_u4_U43 (.A2( u0_u11_u4_n128 ) , .A1( u0_u11_u4_n138 ) , .ZN( u0_u11_u4_n156 ) );
  AOI22_X1 u0_u11_u4_U44 (.B2( u0_u11_u4_n122 ) , .A1( u0_u11_u4_n123 ) , .ZN( u0_u11_u4_n124 ) , .B1( u0_u11_u4_n128 ) , .A2( u0_u11_u4_n172 ) );
  INV_X1 u0_u11_u4_U45 (.A( u0_u11_u4_n153 ) , .ZN( u0_u11_u4_n172 ) );
  NAND2_X1 u0_u11_u4_U46 (.A2( u0_u11_u4_n120 ) , .ZN( u0_u11_u4_n123 ) , .A1( u0_u11_u4_n161 ) );
  AOI22_X1 u0_u11_u4_U47 (.B2( u0_u11_u4_n132 ) , .A2( u0_u11_u4_n133 ) , .ZN( u0_u11_u4_n140 ) , .A1( u0_u11_u4_n150 ) , .B1( u0_u11_u4_n179 ) );
  NAND2_X1 u0_u11_u4_U48 (.ZN( u0_u11_u4_n133 ) , .A2( u0_u11_u4_n146 ) , .A1( u0_u11_u4_n154 ) );
  NAND2_X1 u0_u11_u4_U49 (.A1( u0_u11_u4_n103 ) , .ZN( u0_u11_u4_n154 ) , .A2( u0_u11_u4_n98 ) );
  NOR4_X1 u0_u11_u4_U5 (.A4( u0_u11_u4_n106 ) , .A3( u0_u11_u4_n107 ) , .A2( u0_u11_u4_n108 ) , .A1( u0_u11_u4_n109 ) , .ZN( u0_u11_u4_n110 ) );
  NAND2_X1 u0_u11_u4_U50 (.A1( u0_u11_u4_n101 ) , .ZN( u0_u11_u4_n158 ) , .A2( u0_u11_u4_n99 ) );
  AOI21_X1 u0_u11_u4_U51 (.ZN( u0_u11_u4_n127 ) , .A( u0_u11_u4_n136 ) , .B2( u0_u11_u4_n150 ) , .B1( u0_u11_u4_n180 ) );
  INV_X1 u0_u11_u4_U52 (.A( u0_u11_u4_n160 ) , .ZN( u0_u11_u4_n180 ) );
  NAND2_X1 u0_u11_u4_U53 (.A2( u0_u11_u4_n104 ) , .A1( u0_u11_u4_n105 ) , .ZN( u0_u11_u4_n146 ) );
  NAND2_X1 u0_u11_u4_U54 (.A2( u0_u11_u4_n101 ) , .A1( u0_u11_u4_n102 ) , .ZN( u0_u11_u4_n160 ) );
  NAND2_X1 u0_u11_u4_U55 (.ZN( u0_u11_u4_n134 ) , .A1( u0_u11_u4_n98 ) , .A2( u0_u11_u4_n99 ) );
  NAND2_X1 u0_u11_u4_U56 (.A1( u0_u11_u4_n103 ) , .A2( u0_u11_u4_n104 ) , .ZN( u0_u11_u4_n143 ) );
  NAND2_X1 u0_u11_u4_U57 (.A2( u0_u11_u4_n105 ) , .ZN( u0_u11_u4_n145 ) , .A1( u0_u11_u4_n98 ) );
  NAND2_X1 u0_u11_u4_U58 (.A1( u0_u11_u4_n100 ) , .A2( u0_u11_u4_n105 ) , .ZN( u0_u11_u4_n120 ) );
  NAND2_X1 u0_u11_u4_U59 (.A1( u0_u11_u4_n102 ) , .A2( u0_u11_u4_n104 ) , .ZN( u0_u11_u4_n148 ) );
  AOI21_X1 u0_u11_u4_U6 (.ZN( u0_u11_u4_n106 ) , .B2( u0_u11_u4_n146 ) , .B1( u0_u11_u4_n158 ) , .A( u0_u11_u4_n170 ) );
  NAND2_X1 u0_u11_u4_U60 (.A2( u0_u11_u4_n100 ) , .A1( u0_u11_u4_n103 ) , .ZN( u0_u11_u4_n157 ) );
  INV_X1 u0_u11_u4_U61 (.A( u0_u11_u4_n150 ) , .ZN( u0_u11_u4_n173 ) );
  INV_X1 u0_u11_u4_U62 (.A( u0_u11_u4_n152 ) , .ZN( u0_u11_u4_n171 ) );
  NAND2_X1 u0_u11_u4_U63 (.A1( u0_u11_u4_n100 ) , .ZN( u0_u11_u4_n118 ) , .A2( u0_u11_u4_n99 ) );
  NAND2_X1 u0_u11_u4_U64 (.A2( u0_u11_u4_n100 ) , .A1( u0_u11_u4_n102 ) , .ZN( u0_u11_u4_n144 ) );
  NAND2_X1 u0_u11_u4_U65 (.A2( u0_u11_u4_n101 ) , .A1( u0_u11_u4_n105 ) , .ZN( u0_u11_u4_n96 ) );
  INV_X1 u0_u11_u4_U66 (.A( u0_u11_u4_n128 ) , .ZN( u0_u11_u4_n174 ) );
  NAND2_X1 u0_u11_u4_U67 (.A2( u0_u11_u4_n102 ) , .ZN( u0_u11_u4_n119 ) , .A1( u0_u11_u4_n98 ) );
  NAND2_X1 u0_u11_u4_U68 (.A2( u0_u11_u4_n101 ) , .A1( u0_u11_u4_n103 ) , .ZN( u0_u11_u4_n147 ) );
  NAND2_X1 u0_u11_u4_U69 (.A2( u0_u11_u4_n104 ) , .ZN( u0_u11_u4_n113 ) , .A1( u0_u11_u4_n99 ) );
  AOI21_X1 u0_u11_u4_U7 (.ZN( u0_u11_u4_n108 ) , .B2( u0_u11_u4_n134 ) , .B1( u0_u11_u4_n155 ) , .A( u0_u11_u4_n156 ) );
  NOR2_X1 u0_u11_u4_U70 (.A2( u0_u11_X_28 ) , .ZN( u0_u11_u4_n150 ) , .A1( u0_u11_u4_n168 ) );
  NOR2_X1 u0_u11_u4_U71 (.A2( u0_u11_X_29 ) , .ZN( u0_u11_u4_n152 ) , .A1( u0_u11_u4_n169 ) );
  NOR2_X1 u0_u11_u4_U72 (.A2( u0_u11_X_26 ) , .ZN( u0_u11_u4_n100 ) , .A1( u0_u11_u4_n177 ) );
  NOR2_X1 u0_u11_u4_U73 (.A2( u0_u11_X_30 ) , .ZN( u0_u11_u4_n105 ) , .A1( u0_u11_u4_n176 ) );
  NOR2_X1 u0_u11_u4_U74 (.A2( u0_u11_X_28 ) , .A1( u0_u11_X_29 ) , .ZN( u0_u11_u4_n128 ) );
  NOR2_X1 u0_u11_u4_U75 (.A2( u0_u11_X_25 ) , .A1( u0_u11_X_26 ) , .ZN( u0_u11_u4_n98 ) );
  NOR2_X1 u0_u11_u4_U76 (.A2( u0_u11_X_27 ) , .A1( u0_u11_X_30 ) , .ZN( u0_u11_u4_n102 ) );
  AND2_X1 u0_u11_u4_U77 (.A2( u0_u11_X_25 ) , .A1( u0_u11_X_26 ) , .ZN( u0_u11_u4_n104 ) );
  AND2_X1 u0_u11_u4_U78 (.A1( u0_u11_X_30 ) , .A2( u0_u11_u4_n176 ) , .ZN( u0_u11_u4_n99 ) );
  AND2_X1 u0_u11_u4_U79 (.A1( u0_u11_X_26 ) , .ZN( u0_u11_u4_n101 ) , .A2( u0_u11_u4_n177 ) );
  AOI21_X1 u0_u11_u4_U8 (.ZN( u0_u11_u4_n109 ) , .A( u0_u11_u4_n153 ) , .B1( u0_u11_u4_n159 ) , .B2( u0_u11_u4_n184 ) );
  AND2_X1 u0_u11_u4_U80 (.A1( u0_u11_X_27 ) , .A2( u0_u11_X_30 ) , .ZN( u0_u11_u4_n103 ) );
  INV_X1 u0_u11_u4_U81 (.A( u0_u11_X_28 ) , .ZN( u0_u11_u4_n169 ) );
  INV_X1 u0_u11_u4_U82 (.A( u0_u11_X_29 ) , .ZN( u0_u11_u4_n168 ) );
  INV_X1 u0_u11_u4_U83 (.A( u0_u11_X_25 ) , .ZN( u0_u11_u4_n177 ) );
  INV_X1 u0_u11_u4_U84 (.A( u0_u11_X_27 ) , .ZN( u0_u11_u4_n176 ) );
  NAND4_X1 u0_u11_u4_U85 (.ZN( u0_out11_25 ) , .A4( u0_u11_u4_n139 ) , .A3( u0_u11_u4_n140 ) , .A2( u0_u11_u4_n141 ) , .A1( u0_u11_u4_n142 ) );
  OAI21_X1 u0_u11_u4_U86 (.A( u0_u11_u4_n128 ) , .B2( u0_u11_u4_n129 ) , .B1( u0_u11_u4_n130 ) , .ZN( u0_u11_u4_n142 ) );
  OAI21_X1 u0_u11_u4_U87 (.B2( u0_u11_u4_n131 ) , .ZN( u0_u11_u4_n141 ) , .A( u0_u11_u4_n175 ) , .B1( u0_u11_u4_n183 ) );
  NAND4_X1 u0_u11_u4_U88 (.ZN( u0_out11_14 ) , .A4( u0_u11_u4_n124 ) , .A3( u0_u11_u4_n125 ) , .A2( u0_u11_u4_n126 ) , .A1( u0_u11_u4_n127 ) );
  AOI22_X1 u0_u11_u4_U89 (.B2( u0_u11_u4_n117 ) , .ZN( u0_u11_u4_n126 ) , .A1( u0_u11_u4_n129 ) , .B1( u0_u11_u4_n152 ) , .A2( u0_u11_u4_n175 ) );
  AOI211_X1 u0_u11_u4_U9 (.B( u0_u11_u4_n136 ) , .A( u0_u11_u4_n137 ) , .C2( u0_u11_u4_n138 ) , .ZN( u0_u11_u4_n139 ) , .C1( u0_u11_u4_n182 ) );
  AOI22_X1 u0_u11_u4_U90 (.ZN( u0_u11_u4_n125 ) , .B2( u0_u11_u4_n131 ) , .A2( u0_u11_u4_n132 ) , .B1( u0_u11_u4_n138 ) , .A1( u0_u11_u4_n178 ) );
  NAND4_X1 u0_u11_u4_U91 (.ZN( u0_out11_8 ) , .A4( u0_u11_u4_n110 ) , .A3( u0_u11_u4_n111 ) , .A2( u0_u11_u4_n112 ) , .A1( u0_u11_u4_n186 ) );
  NAND2_X1 u0_u11_u4_U92 (.ZN( u0_u11_u4_n112 ) , .A2( u0_u11_u4_n130 ) , .A1( u0_u11_u4_n150 ) );
  AOI22_X1 u0_u11_u4_U93 (.ZN( u0_u11_u4_n111 ) , .B2( u0_u11_u4_n132 ) , .A1( u0_u11_u4_n152 ) , .B1( u0_u11_u4_n178 ) , .A2( u0_u11_u4_n97 ) );
  AOI22_X1 u0_u11_u4_U94 (.B2( u0_u11_u4_n149 ) , .B1( u0_u11_u4_n150 ) , .A2( u0_u11_u4_n151 ) , .A1( u0_u11_u4_n152 ) , .ZN( u0_u11_u4_n167 ) );
  NOR4_X1 u0_u11_u4_U95 (.A4( u0_u11_u4_n162 ) , .A3( u0_u11_u4_n163 ) , .A2( u0_u11_u4_n164 ) , .A1( u0_u11_u4_n165 ) , .ZN( u0_u11_u4_n166 ) );
  NAND3_X1 u0_u11_u4_U96 (.ZN( u0_out11_3 ) , .A3( u0_u11_u4_n166 ) , .A1( u0_u11_u4_n167 ) , .A2( u0_u11_u4_n186 ) );
  NAND3_X1 u0_u11_u4_U97 (.A3( u0_u11_u4_n146 ) , .A2( u0_u11_u4_n147 ) , .A1( u0_u11_u4_n148 ) , .ZN( u0_u11_u4_n149 ) );
  NAND3_X1 u0_u11_u4_U98 (.A3( u0_u11_u4_n143 ) , .A2( u0_u11_u4_n144 ) , .A1( u0_u11_u4_n145 ) , .ZN( u0_u11_u4_n151 ) );
  NAND3_X1 u0_u11_u4_U99 (.A3( u0_u11_u4_n121 ) , .ZN( u0_u11_u4_n122 ) , .A2( u0_u11_u4_n144 ) , .A1( u0_u11_u4_n154 ) );
  INV_X1 u0_u11_u5_U10 (.A( u0_u11_u5_n121 ) , .ZN( u0_u11_u5_n177 ) );
  NOR3_X1 u0_u11_u5_U100 (.A3( u0_u11_u5_n141 ) , .A1( u0_u11_u5_n142 ) , .ZN( u0_u11_u5_n143 ) , .A2( u0_u11_u5_n191 ) );
  NAND4_X1 u0_u11_u5_U101 (.ZN( u0_out11_4 ) , .A4( u0_u11_u5_n112 ) , .A2( u0_u11_u5_n113 ) , .A1( u0_u11_u5_n114 ) , .A3( u0_u11_u5_n195 ) );
  AOI211_X1 u0_u11_u5_U102 (.A( u0_u11_u5_n110 ) , .C1( u0_u11_u5_n111 ) , .ZN( u0_u11_u5_n112 ) , .B( u0_u11_u5_n118 ) , .C2( u0_u11_u5_n177 ) );
  AOI222_X1 u0_u11_u5_U103 (.ZN( u0_u11_u5_n113 ) , .A1( u0_u11_u5_n131 ) , .C1( u0_u11_u5_n148 ) , .B2( u0_u11_u5_n174 ) , .C2( u0_u11_u5_n178 ) , .A2( u0_u11_u5_n179 ) , .B1( u0_u11_u5_n99 ) );
  NAND3_X1 u0_u11_u5_U104 (.A2( u0_u11_u5_n154 ) , .A3( u0_u11_u5_n158 ) , .A1( u0_u11_u5_n161 ) , .ZN( u0_u11_u5_n99 ) );
  NOR2_X1 u0_u11_u5_U11 (.ZN( u0_u11_u5_n160 ) , .A2( u0_u11_u5_n173 ) , .A1( u0_u11_u5_n177 ) );
  INV_X1 u0_u11_u5_U12 (.A( u0_u11_u5_n150 ) , .ZN( u0_u11_u5_n174 ) );
  AOI21_X1 u0_u11_u5_U13 (.A( u0_u11_u5_n160 ) , .B2( u0_u11_u5_n161 ) , .ZN( u0_u11_u5_n162 ) , .B1( u0_u11_u5_n192 ) );
  INV_X1 u0_u11_u5_U14 (.A( u0_u11_u5_n159 ) , .ZN( u0_u11_u5_n192 ) );
  AOI21_X1 u0_u11_u5_U15 (.A( u0_u11_u5_n156 ) , .B2( u0_u11_u5_n157 ) , .B1( u0_u11_u5_n158 ) , .ZN( u0_u11_u5_n163 ) );
  AOI21_X1 u0_u11_u5_U16 (.B2( u0_u11_u5_n139 ) , .B1( u0_u11_u5_n140 ) , .ZN( u0_u11_u5_n141 ) , .A( u0_u11_u5_n150 ) );
  OAI21_X1 u0_u11_u5_U17 (.A( u0_u11_u5_n133 ) , .B2( u0_u11_u5_n134 ) , .B1( u0_u11_u5_n135 ) , .ZN( u0_u11_u5_n142 ) );
  OAI21_X1 u0_u11_u5_U18 (.ZN( u0_u11_u5_n133 ) , .B2( u0_u11_u5_n147 ) , .A( u0_u11_u5_n173 ) , .B1( u0_u11_u5_n188 ) );
  NAND2_X1 u0_u11_u5_U19 (.A2( u0_u11_u5_n119 ) , .A1( u0_u11_u5_n123 ) , .ZN( u0_u11_u5_n137 ) );
  INV_X1 u0_u11_u5_U20 (.A( u0_u11_u5_n155 ) , .ZN( u0_u11_u5_n194 ) );
  NAND2_X1 u0_u11_u5_U21 (.A1( u0_u11_u5_n121 ) , .ZN( u0_u11_u5_n132 ) , .A2( u0_u11_u5_n172 ) );
  NAND2_X1 u0_u11_u5_U22 (.A2( u0_u11_u5_n122 ) , .ZN( u0_u11_u5_n136 ) , .A1( u0_u11_u5_n154 ) );
  NAND2_X1 u0_u11_u5_U23 (.A2( u0_u11_u5_n119 ) , .A1( u0_u11_u5_n120 ) , .ZN( u0_u11_u5_n159 ) );
  INV_X1 u0_u11_u5_U24 (.A( u0_u11_u5_n156 ) , .ZN( u0_u11_u5_n175 ) );
  INV_X1 u0_u11_u5_U25 (.A( u0_u11_u5_n158 ) , .ZN( u0_u11_u5_n188 ) );
  INV_X1 u0_u11_u5_U26 (.A( u0_u11_u5_n152 ) , .ZN( u0_u11_u5_n179 ) );
  INV_X1 u0_u11_u5_U27 (.A( u0_u11_u5_n140 ) , .ZN( u0_u11_u5_n182 ) );
  INV_X1 u0_u11_u5_U28 (.A( u0_u11_u5_n151 ) , .ZN( u0_u11_u5_n183 ) );
  INV_X1 u0_u11_u5_U29 (.A( u0_u11_u5_n123 ) , .ZN( u0_u11_u5_n185 ) );
  NOR2_X1 u0_u11_u5_U3 (.ZN( u0_u11_u5_n134 ) , .A1( u0_u11_u5_n183 ) , .A2( u0_u11_u5_n190 ) );
  INV_X1 u0_u11_u5_U30 (.A( u0_u11_u5_n161 ) , .ZN( u0_u11_u5_n184 ) );
  INV_X1 u0_u11_u5_U31 (.A( u0_u11_u5_n139 ) , .ZN( u0_u11_u5_n189 ) );
  INV_X1 u0_u11_u5_U32 (.A( u0_u11_u5_n157 ) , .ZN( u0_u11_u5_n190 ) );
  INV_X1 u0_u11_u5_U33 (.A( u0_u11_u5_n120 ) , .ZN( u0_u11_u5_n193 ) );
  NAND2_X1 u0_u11_u5_U34 (.ZN( u0_u11_u5_n111 ) , .A1( u0_u11_u5_n140 ) , .A2( u0_u11_u5_n155 ) );
  NOR2_X1 u0_u11_u5_U35 (.ZN( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n170 ) , .A2( u0_u11_u5_n180 ) );
  INV_X1 u0_u11_u5_U36 (.A( u0_u11_u5_n117 ) , .ZN( u0_u11_u5_n196 ) );
  OAI221_X1 u0_u11_u5_U37 (.A( u0_u11_u5_n116 ) , .ZN( u0_u11_u5_n117 ) , .B2( u0_u11_u5_n119 ) , .C1( u0_u11_u5_n153 ) , .C2( u0_u11_u5_n158 ) , .B1( u0_u11_u5_n172 ) );
  AOI222_X1 u0_u11_u5_U38 (.ZN( u0_u11_u5_n116 ) , .B2( u0_u11_u5_n145 ) , .C1( u0_u11_u5_n148 ) , .A2( u0_u11_u5_n174 ) , .C2( u0_u11_u5_n177 ) , .B1( u0_u11_u5_n187 ) , .A1( u0_u11_u5_n193 ) );
  INV_X1 u0_u11_u5_U39 (.A( u0_u11_u5_n115 ) , .ZN( u0_u11_u5_n187 ) );
  INV_X1 u0_u11_u5_U4 (.A( u0_u11_u5_n138 ) , .ZN( u0_u11_u5_n191 ) );
  AOI22_X1 u0_u11_u5_U40 (.B2( u0_u11_u5_n131 ) , .A2( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n169 ) , .B1( u0_u11_u5_n174 ) , .A1( u0_u11_u5_n185 ) );
  NOR2_X1 u0_u11_u5_U41 (.A1( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n150 ) , .A2( u0_u11_u5_n173 ) );
  AOI21_X1 u0_u11_u5_U42 (.A( u0_u11_u5_n118 ) , .B2( u0_u11_u5_n145 ) , .ZN( u0_u11_u5_n168 ) , .B1( u0_u11_u5_n186 ) );
  INV_X1 u0_u11_u5_U43 (.A( u0_u11_u5_n122 ) , .ZN( u0_u11_u5_n186 ) );
  NOR2_X1 u0_u11_u5_U44 (.A1( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n152 ) , .A2( u0_u11_u5_n176 ) );
  NOR2_X1 u0_u11_u5_U45 (.A1( u0_u11_u5_n115 ) , .ZN( u0_u11_u5_n118 ) , .A2( u0_u11_u5_n153 ) );
  NOR2_X1 u0_u11_u5_U46 (.A2( u0_u11_u5_n145 ) , .ZN( u0_u11_u5_n156 ) , .A1( u0_u11_u5_n174 ) );
  NOR2_X1 u0_u11_u5_U47 (.ZN( u0_u11_u5_n121 ) , .A2( u0_u11_u5_n145 ) , .A1( u0_u11_u5_n176 ) );
  AOI22_X1 u0_u11_u5_U48 (.ZN( u0_u11_u5_n114 ) , .A2( u0_u11_u5_n137 ) , .A1( u0_u11_u5_n145 ) , .B2( u0_u11_u5_n175 ) , .B1( u0_u11_u5_n193 ) );
  OAI211_X1 u0_u11_u5_U49 (.B( u0_u11_u5_n124 ) , .A( u0_u11_u5_n125 ) , .C2( u0_u11_u5_n126 ) , .C1( u0_u11_u5_n127 ) , .ZN( u0_u11_u5_n128 ) );
  OAI21_X1 u0_u11_u5_U5 (.B2( u0_u11_u5_n136 ) , .B1( u0_u11_u5_n137 ) , .ZN( u0_u11_u5_n138 ) , .A( u0_u11_u5_n177 ) );
  OAI21_X1 u0_u11_u5_U50 (.ZN( u0_u11_u5_n124 ) , .A( u0_u11_u5_n177 ) , .B2( u0_u11_u5_n183 ) , .B1( u0_u11_u5_n189 ) );
  NOR3_X1 u0_u11_u5_U51 (.ZN( u0_u11_u5_n127 ) , .A1( u0_u11_u5_n136 ) , .A3( u0_u11_u5_n148 ) , .A2( u0_u11_u5_n182 ) );
  OAI21_X1 u0_u11_u5_U52 (.ZN( u0_u11_u5_n125 ) , .A( u0_u11_u5_n174 ) , .B2( u0_u11_u5_n185 ) , .B1( u0_u11_u5_n190 ) );
  AOI21_X1 u0_u11_u5_U53 (.A( u0_u11_u5_n153 ) , .B2( u0_u11_u5_n154 ) , .B1( u0_u11_u5_n155 ) , .ZN( u0_u11_u5_n164 ) );
  AOI21_X1 u0_u11_u5_U54 (.ZN( u0_u11_u5_n110 ) , .B1( u0_u11_u5_n122 ) , .B2( u0_u11_u5_n139 ) , .A( u0_u11_u5_n153 ) );
  INV_X1 u0_u11_u5_U55 (.A( u0_u11_u5_n153 ) , .ZN( u0_u11_u5_n176 ) );
  INV_X1 u0_u11_u5_U56 (.A( u0_u11_u5_n126 ) , .ZN( u0_u11_u5_n173 ) );
  AND2_X1 u0_u11_u5_U57 (.A2( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n107 ) , .ZN( u0_u11_u5_n147 ) );
  AND2_X1 u0_u11_u5_U58 (.A2( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n108 ) , .ZN( u0_u11_u5_n148 ) );
  NAND2_X1 u0_u11_u5_U59 (.A1( u0_u11_u5_n105 ) , .A2( u0_u11_u5_n106 ) , .ZN( u0_u11_u5_n158 ) );
  INV_X1 u0_u11_u5_U6 (.A( u0_u11_u5_n135 ) , .ZN( u0_u11_u5_n178 ) );
  NAND2_X1 u0_u11_u5_U60 (.A2( u0_u11_u5_n108 ) , .A1( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n139 ) );
  NAND2_X1 u0_u11_u5_U61 (.A1( u0_u11_u5_n106 ) , .A2( u0_u11_u5_n108 ) , .ZN( u0_u11_u5_n119 ) );
  NAND2_X1 u0_u11_u5_U62 (.A2( u0_u11_u5_n103 ) , .A1( u0_u11_u5_n105 ) , .ZN( u0_u11_u5_n140 ) );
  NAND2_X1 u0_u11_u5_U63 (.A2( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n105 ) , .ZN( u0_u11_u5_n155 ) );
  NAND2_X1 u0_u11_u5_U64 (.A2( u0_u11_u5_n106 ) , .A1( u0_u11_u5_n107 ) , .ZN( u0_u11_u5_n122 ) );
  NAND2_X1 u0_u11_u5_U65 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n106 ) , .ZN( u0_u11_u5_n115 ) );
  NAND2_X1 u0_u11_u5_U66 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n103 ) , .ZN( u0_u11_u5_n161 ) );
  NAND2_X1 u0_u11_u5_U67 (.A1( u0_u11_u5_n105 ) , .A2( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n154 ) );
  INV_X1 u0_u11_u5_U68 (.A( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n172 ) );
  NAND2_X1 u0_u11_u5_U69 (.A1( u0_u11_u5_n103 ) , .A2( u0_u11_u5_n108 ) , .ZN( u0_u11_u5_n123 ) );
  OAI22_X1 u0_u11_u5_U7 (.B2( u0_u11_u5_n149 ) , .B1( u0_u11_u5_n150 ) , .A2( u0_u11_u5_n151 ) , .A1( u0_u11_u5_n152 ) , .ZN( u0_u11_u5_n165 ) );
  NAND2_X1 u0_u11_u5_U70 (.A2( u0_u11_u5_n103 ) , .A1( u0_u11_u5_n107 ) , .ZN( u0_u11_u5_n151 ) );
  NAND2_X1 u0_u11_u5_U71 (.A2( u0_u11_u5_n107 ) , .A1( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n120 ) );
  NAND2_X1 u0_u11_u5_U72 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n109 ) , .ZN( u0_u11_u5_n157 ) );
  AND2_X1 u0_u11_u5_U73 (.A2( u0_u11_u5_n100 ) , .A1( u0_u11_u5_n104 ) , .ZN( u0_u11_u5_n131 ) );
  INV_X1 u0_u11_u5_U74 (.A( u0_u11_u5_n102 ) , .ZN( u0_u11_u5_n195 ) );
  OAI221_X1 u0_u11_u5_U75 (.A( u0_u11_u5_n101 ) , .ZN( u0_u11_u5_n102 ) , .C2( u0_u11_u5_n115 ) , .C1( u0_u11_u5_n126 ) , .B1( u0_u11_u5_n134 ) , .B2( u0_u11_u5_n160 ) );
  OAI21_X1 u0_u11_u5_U76 (.ZN( u0_u11_u5_n101 ) , .B1( u0_u11_u5_n137 ) , .A( u0_u11_u5_n146 ) , .B2( u0_u11_u5_n147 ) );
  NOR2_X1 u0_u11_u5_U77 (.A2( u0_u11_X_34 ) , .A1( u0_u11_X_35 ) , .ZN( u0_u11_u5_n145 ) );
  NOR2_X1 u0_u11_u5_U78 (.A2( u0_u11_X_34 ) , .ZN( u0_u11_u5_n146 ) , .A1( u0_u11_u5_n171 ) );
  NOR2_X1 u0_u11_u5_U79 (.A2( u0_u11_X_31 ) , .A1( u0_u11_X_32 ) , .ZN( u0_u11_u5_n103 ) );
  NOR3_X1 u0_u11_u5_U8 (.A2( u0_u11_u5_n147 ) , .A1( u0_u11_u5_n148 ) , .ZN( u0_u11_u5_n149 ) , .A3( u0_u11_u5_n194 ) );
  NOR2_X1 u0_u11_u5_U80 (.A2( u0_u11_X_36 ) , .ZN( u0_u11_u5_n105 ) , .A1( u0_u11_u5_n180 ) );
  NOR2_X1 u0_u11_u5_U81 (.A2( u0_u11_X_33 ) , .ZN( u0_u11_u5_n108 ) , .A1( u0_u11_u5_n170 ) );
  NOR2_X1 u0_u11_u5_U82 (.A2( u0_u11_X_33 ) , .A1( u0_u11_X_36 ) , .ZN( u0_u11_u5_n107 ) );
  NOR2_X1 u0_u11_u5_U83 (.A2( u0_u11_X_31 ) , .ZN( u0_u11_u5_n104 ) , .A1( u0_u11_u5_n181 ) );
  NAND2_X1 u0_u11_u5_U84 (.A2( u0_u11_X_34 ) , .A1( u0_u11_X_35 ) , .ZN( u0_u11_u5_n153 ) );
  NAND2_X1 u0_u11_u5_U85 (.A1( u0_u11_X_34 ) , .ZN( u0_u11_u5_n126 ) , .A2( u0_u11_u5_n171 ) );
  AND2_X1 u0_u11_u5_U86 (.A1( u0_u11_X_31 ) , .A2( u0_u11_X_32 ) , .ZN( u0_u11_u5_n106 ) );
  AND2_X1 u0_u11_u5_U87 (.A1( u0_u11_X_31 ) , .ZN( u0_u11_u5_n109 ) , .A2( u0_u11_u5_n181 ) );
  INV_X1 u0_u11_u5_U88 (.A( u0_u11_X_33 ) , .ZN( u0_u11_u5_n180 ) );
  INV_X1 u0_u11_u5_U89 (.A( u0_u11_X_35 ) , .ZN( u0_u11_u5_n171 ) );
  NOR2_X1 u0_u11_u5_U9 (.ZN( u0_u11_u5_n135 ) , .A1( u0_u11_u5_n173 ) , .A2( u0_u11_u5_n176 ) );
  INV_X1 u0_u11_u5_U90 (.A( u0_u11_X_36 ) , .ZN( u0_u11_u5_n170 ) );
  INV_X1 u0_u11_u5_U91 (.A( u0_u11_X_32 ) , .ZN( u0_u11_u5_n181 ) );
  NAND4_X1 u0_u11_u5_U92 (.ZN( u0_out11_29 ) , .A4( u0_u11_u5_n129 ) , .A3( u0_u11_u5_n130 ) , .A2( u0_u11_u5_n168 ) , .A1( u0_u11_u5_n196 ) );
  AOI221_X1 u0_u11_u5_U93 (.A( u0_u11_u5_n128 ) , .ZN( u0_u11_u5_n129 ) , .C2( u0_u11_u5_n132 ) , .B2( u0_u11_u5_n159 ) , .B1( u0_u11_u5_n176 ) , .C1( u0_u11_u5_n184 ) );
  AOI222_X1 u0_u11_u5_U94 (.ZN( u0_u11_u5_n130 ) , .A2( u0_u11_u5_n146 ) , .B1( u0_u11_u5_n147 ) , .C2( u0_u11_u5_n175 ) , .B2( u0_u11_u5_n179 ) , .A1( u0_u11_u5_n188 ) , .C1( u0_u11_u5_n194 ) );
  NAND4_X1 u0_u11_u5_U95 (.ZN( u0_out11_19 ) , .A4( u0_u11_u5_n166 ) , .A3( u0_u11_u5_n167 ) , .A2( u0_u11_u5_n168 ) , .A1( u0_u11_u5_n169 ) );
  AOI22_X1 u0_u11_u5_U96 (.B2( u0_u11_u5_n145 ) , .A2( u0_u11_u5_n146 ) , .ZN( u0_u11_u5_n167 ) , .B1( u0_u11_u5_n182 ) , .A1( u0_u11_u5_n189 ) );
  NOR4_X1 u0_u11_u5_U97 (.A4( u0_u11_u5_n162 ) , .A3( u0_u11_u5_n163 ) , .A2( u0_u11_u5_n164 ) , .A1( u0_u11_u5_n165 ) , .ZN( u0_u11_u5_n166 ) );
  NAND4_X1 u0_u11_u5_U98 (.ZN( u0_out11_11 ) , .A4( u0_u11_u5_n143 ) , .A3( u0_u11_u5_n144 ) , .A2( u0_u11_u5_n169 ) , .A1( u0_u11_u5_n196 ) );
  AOI22_X1 u0_u11_u5_U99 (.A2( u0_u11_u5_n132 ) , .ZN( u0_u11_u5_n144 ) , .B2( u0_u11_u5_n145 ) , .B1( u0_u11_u5_n184 ) , .A1( u0_u11_u5_n194 ) );
  OAI21_X1 u0_u11_u6_U10 (.A( u0_u11_u6_n159 ) , .B1( u0_u11_u6_n169 ) , .B2( u0_u11_u6_n173 ) , .ZN( u0_u11_u6_n90 ) );
  INV_X1 u0_u11_u6_U11 (.ZN( u0_u11_u6_n172 ) , .A( u0_u11_u6_n88 ) );
  AOI22_X1 u0_u11_u6_U12 (.A2( u0_u11_u6_n151 ) , .B2( u0_u11_u6_n161 ) , .A1( u0_u11_u6_n167 ) , .B1( u0_u11_u6_n170 ) , .ZN( u0_u11_u6_n89 ) );
  AOI21_X1 u0_u11_u6_U13 (.ZN( u0_u11_u6_n106 ) , .A( u0_u11_u6_n142 ) , .B2( u0_u11_u6_n159 ) , .B1( u0_u11_u6_n164 ) );
  INV_X1 u0_u11_u6_U14 (.A( u0_u11_u6_n155 ) , .ZN( u0_u11_u6_n161 ) );
  INV_X1 u0_u11_u6_U15 (.A( u0_u11_u6_n128 ) , .ZN( u0_u11_u6_n164 ) );
  NAND2_X1 u0_u11_u6_U16 (.ZN( u0_u11_u6_n110 ) , .A1( u0_u11_u6_n122 ) , .A2( u0_u11_u6_n129 ) );
  NAND2_X1 u0_u11_u6_U17 (.ZN( u0_u11_u6_n124 ) , .A2( u0_u11_u6_n146 ) , .A1( u0_u11_u6_n148 ) );
  INV_X1 u0_u11_u6_U18 (.A( u0_u11_u6_n132 ) , .ZN( u0_u11_u6_n171 ) );
  AND2_X1 u0_u11_u6_U19 (.A1( u0_u11_u6_n100 ) , .ZN( u0_u11_u6_n130 ) , .A2( u0_u11_u6_n147 ) );
  INV_X1 u0_u11_u6_U20 (.A( u0_u11_u6_n127 ) , .ZN( u0_u11_u6_n173 ) );
  INV_X1 u0_u11_u6_U21 (.A( u0_u11_u6_n121 ) , .ZN( u0_u11_u6_n167 ) );
  INV_X1 u0_u11_u6_U22 (.A( u0_u11_u6_n100 ) , .ZN( u0_u11_u6_n169 ) );
  INV_X1 u0_u11_u6_U23 (.A( u0_u11_u6_n123 ) , .ZN( u0_u11_u6_n170 ) );
  INV_X1 u0_u11_u6_U24 (.A( u0_u11_u6_n113 ) , .ZN( u0_u11_u6_n168 ) );
  AND2_X1 u0_u11_u6_U25 (.A1( u0_u11_u6_n107 ) , .A2( u0_u11_u6_n119 ) , .ZN( u0_u11_u6_n133 ) );
  AND2_X1 u0_u11_u6_U26 (.A2( u0_u11_u6_n121 ) , .A1( u0_u11_u6_n122 ) , .ZN( u0_u11_u6_n131 ) );
  AND3_X1 u0_u11_u6_U27 (.ZN( u0_u11_u6_n120 ) , .A2( u0_u11_u6_n127 ) , .A1( u0_u11_u6_n132 ) , .A3( u0_u11_u6_n145 ) );
  INV_X1 u0_u11_u6_U28 (.A( u0_u11_u6_n146 ) , .ZN( u0_u11_u6_n163 ) );
  AOI222_X1 u0_u11_u6_U29 (.ZN( u0_u11_u6_n114 ) , .A1( u0_u11_u6_n118 ) , .A2( u0_u11_u6_n126 ) , .B2( u0_u11_u6_n151 ) , .C2( u0_u11_u6_n159 ) , .C1( u0_u11_u6_n168 ) , .B1( u0_u11_u6_n169 ) );
  INV_X1 u0_u11_u6_U3 (.A( u0_u11_u6_n110 ) , .ZN( u0_u11_u6_n166 ) );
  NOR2_X1 u0_u11_u6_U30 (.A1( u0_u11_u6_n162 ) , .A2( u0_u11_u6_n165 ) , .ZN( u0_u11_u6_n98 ) );
  NAND2_X1 u0_u11_u6_U31 (.A1( u0_u11_u6_n144 ) , .ZN( u0_u11_u6_n151 ) , .A2( u0_u11_u6_n158 ) );
  NAND2_X1 u0_u11_u6_U32 (.ZN( u0_u11_u6_n132 ) , .A1( u0_u11_u6_n91 ) , .A2( u0_u11_u6_n97 ) );
  AOI22_X1 u0_u11_u6_U33 (.B2( u0_u11_u6_n110 ) , .B1( u0_u11_u6_n111 ) , .A1( u0_u11_u6_n112 ) , .ZN( u0_u11_u6_n115 ) , .A2( u0_u11_u6_n161 ) );
  NAND4_X1 u0_u11_u6_U34 (.A3( u0_u11_u6_n109 ) , .ZN( u0_u11_u6_n112 ) , .A4( u0_u11_u6_n132 ) , .A2( u0_u11_u6_n147 ) , .A1( u0_u11_u6_n166 ) );
  NOR2_X1 u0_u11_u6_U35 (.ZN( u0_u11_u6_n109 ) , .A1( u0_u11_u6_n170 ) , .A2( u0_u11_u6_n173 ) );
  NOR2_X1 u0_u11_u6_U36 (.A2( u0_u11_u6_n126 ) , .ZN( u0_u11_u6_n155 ) , .A1( u0_u11_u6_n160 ) );
  NAND2_X1 u0_u11_u6_U37 (.ZN( u0_u11_u6_n146 ) , .A2( u0_u11_u6_n94 ) , .A1( u0_u11_u6_n99 ) );
  AOI21_X1 u0_u11_u6_U38 (.A( u0_u11_u6_n144 ) , .B2( u0_u11_u6_n145 ) , .B1( u0_u11_u6_n146 ) , .ZN( u0_u11_u6_n150 ) );
  AOI211_X1 u0_u11_u6_U39 (.B( u0_u11_u6_n134 ) , .A( u0_u11_u6_n135 ) , .C1( u0_u11_u6_n136 ) , .ZN( u0_u11_u6_n137 ) , .C2( u0_u11_u6_n151 ) );
  INV_X1 u0_u11_u6_U4 (.A( u0_u11_u6_n142 ) , .ZN( u0_u11_u6_n174 ) );
  NAND4_X1 u0_u11_u6_U40 (.A4( u0_u11_u6_n127 ) , .A3( u0_u11_u6_n128 ) , .A2( u0_u11_u6_n129 ) , .A1( u0_u11_u6_n130 ) , .ZN( u0_u11_u6_n136 ) );
  AOI21_X1 u0_u11_u6_U41 (.B2( u0_u11_u6_n132 ) , .B1( u0_u11_u6_n133 ) , .ZN( u0_u11_u6_n134 ) , .A( u0_u11_u6_n158 ) );
  AOI21_X1 u0_u11_u6_U42 (.B1( u0_u11_u6_n131 ) , .ZN( u0_u11_u6_n135 ) , .A( u0_u11_u6_n144 ) , .B2( u0_u11_u6_n146 ) );
  INV_X1 u0_u11_u6_U43 (.A( u0_u11_u6_n111 ) , .ZN( u0_u11_u6_n158 ) );
  NAND2_X1 u0_u11_u6_U44 (.ZN( u0_u11_u6_n127 ) , .A1( u0_u11_u6_n91 ) , .A2( u0_u11_u6_n92 ) );
  NAND2_X1 u0_u11_u6_U45 (.ZN( u0_u11_u6_n129 ) , .A2( u0_u11_u6_n95 ) , .A1( u0_u11_u6_n96 ) );
  INV_X1 u0_u11_u6_U46 (.A( u0_u11_u6_n144 ) , .ZN( u0_u11_u6_n159 ) );
  NAND2_X1 u0_u11_u6_U47 (.ZN( u0_u11_u6_n145 ) , .A2( u0_u11_u6_n97 ) , .A1( u0_u11_u6_n98 ) );
  NAND2_X1 u0_u11_u6_U48 (.ZN( u0_u11_u6_n148 ) , .A2( u0_u11_u6_n92 ) , .A1( u0_u11_u6_n94 ) );
  NAND2_X1 u0_u11_u6_U49 (.ZN( u0_u11_u6_n108 ) , .A2( u0_u11_u6_n139 ) , .A1( u0_u11_u6_n144 ) );
  NAND2_X1 u0_u11_u6_U5 (.A2( u0_u11_u6_n143 ) , .ZN( u0_u11_u6_n152 ) , .A1( u0_u11_u6_n166 ) );
  NAND2_X1 u0_u11_u6_U50 (.ZN( u0_u11_u6_n121 ) , .A2( u0_u11_u6_n95 ) , .A1( u0_u11_u6_n97 ) );
  NAND2_X1 u0_u11_u6_U51 (.ZN( u0_u11_u6_n107 ) , .A2( u0_u11_u6_n92 ) , .A1( u0_u11_u6_n95 ) );
  AND2_X1 u0_u11_u6_U52 (.ZN( u0_u11_u6_n118 ) , .A2( u0_u11_u6_n91 ) , .A1( u0_u11_u6_n99 ) );
  NAND2_X1 u0_u11_u6_U53 (.ZN( u0_u11_u6_n147 ) , .A2( u0_u11_u6_n98 ) , .A1( u0_u11_u6_n99 ) );
  NAND2_X1 u0_u11_u6_U54 (.ZN( u0_u11_u6_n128 ) , .A1( u0_u11_u6_n94 ) , .A2( u0_u11_u6_n96 ) );
  NAND2_X1 u0_u11_u6_U55 (.ZN( u0_u11_u6_n119 ) , .A2( u0_u11_u6_n95 ) , .A1( u0_u11_u6_n99 ) );
  NAND2_X1 u0_u11_u6_U56 (.ZN( u0_u11_u6_n123 ) , .A2( u0_u11_u6_n91 ) , .A1( u0_u11_u6_n96 ) );
  NAND2_X1 u0_u11_u6_U57 (.ZN( u0_u11_u6_n100 ) , .A2( u0_u11_u6_n92 ) , .A1( u0_u11_u6_n98 ) );
  NAND2_X1 u0_u11_u6_U58 (.ZN( u0_u11_u6_n122 ) , .A1( u0_u11_u6_n94 ) , .A2( u0_u11_u6_n97 ) );
  INV_X1 u0_u11_u6_U59 (.A( u0_u11_u6_n139 ) , .ZN( u0_u11_u6_n160 ) );
  AOI22_X1 u0_u11_u6_U6 (.B2( u0_u11_u6_n101 ) , .A1( u0_u11_u6_n102 ) , .ZN( u0_u11_u6_n103 ) , .B1( u0_u11_u6_n160 ) , .A2( u0_u11_u6_n161 ) );
  NAND2_X1 u0_u11_u6_U60 (.ZN( u0_u11_u6_n113 ) , .A1( u0_u11_u6_n96 ) , .A2( u0_u11_u6_n98 ) );
  NOR2_X1 u0_u11_u6_U61 (.A2( u0_u11_X_40 ) , .A1( u0_u11_X_41 ) , .ZN( u0_u11_u6_n126 ) );
  NOR2_X1 u0_u11_u6_U62 (.A2( u0_u11_X_39 ) , .A1( u0_u11_X_42 ) , .ZN( u0_u11_u6_n92 ) );
  NOR2_X1 u0_u11_u6_U63 (.A2( u0_u11_X_39 ) , .A1( u0_u11_u6_n156 ) , .ZN( u0_u11_u6_n97 ) );
  NOR2_X1 u0_u11_u6_U64 (.A2( u0_u11_X_38 ) , .A1( u0_u11_u6_n165 ) , .ZN( u0_u11_u6_n95 ) );
  NOR2_X1 u0_u11_u6_U65 (.A2( u0_u11_X_41 ) , .ZN( u0_u11_u6_n111 ) , .A1( u0_u11_u6_n157 ) );
  NOR2_X1 u0_u11_u6_U66 (.A2( u0_u11_X_37 ) , .A1( u0_u11_u6_n162 ) , .ZN( u0_u11_u6_n94 ) );
  NOR2_X1 u0_u11_u6_U67 (.A2( u0_u11_X_37 ) , .A1( u0_u11_X_38 ) , .ZN( u0_u11_u6_n91 ) );
  NAND2_X1 u0_u11_u6_U68 (.A1( u0_u11_X_41 ) , .ZN( u0_u11_u6_n144 ) , .A2( u0_u11_u6_n157 ) );
  NAND2_X1 u0_u11_u6_U69 (.A2( u0_u11_X_40 ) , .A1( u0_u11_X_41 ) , .ZN( u0_u11_u6_n139 ) );
  NOR2_X1 u0_u11_u6_U7 (.A1( u0_u11_u6_n118 ) , .ZN( u0_u11_u6_n143 ) , .A2( u0_u11_u6_n168 ) );
  AND2_X1 u0_u11_u6_U70 (.A1( u0_u11_X_39 ) , .A2( u0_u11_u6_n156 ) , .ZN( u0_u11_u6_n96 ) );
  AND2_X1 u0_u11_u6_U71 (.A1( u0_u11_X_39 ) , .A2( u0_u11_X_42 ) , .ZN( u0_u11_u6_n99 ) );
  INV_X1 u0_u11_u6_U72 (.A( u0_u11_X_40 ) , .ZN( u0_u11_u6_n157 ) );
  INV_X1 u0_u11_u6_U73 (.A( u0_u11_X_37 ) , .ZN( u0_u11_u6_n165 ) );
  INV_X1 u0_u11_u6_U74 (.A( u0_u11_X_38 ) , .ZN( u0_u11_u6_n162 ) );
  INV_X1 u0_u11_u6_U75 (.A( u0_u11_X_42 ) , .ZN( u0_u11_u6_n156 ) );
  NAND4_X1 u0_u11_u6_U76 (.ZN( u0_out11_32 ) , .A4( u0_u11_u6_n103 ) , .A3( u0_u11_u6_n104 ) , .A2( u0_u11_u6_n105 ) , .A1( u0_u11_u6_n106 ) );
  AOI22_X1 u0_u11_u6_U77 (.ZN( u0_u11_u6_n105 ) , .A2( u0_u11_u6_n108 ) , .A1( u0_u11_u6_n118 ) , .B2( u0_u11_u6_n126 ) , .B1( u0_u11_u6_n171 ) );
  AOI22_X1 u0_u11_u6_U78 (.ZN( u0_u11_u6_n104 ) , .A1( u0_u11_u6_n111 ) , .B1( u0_u11_u6_n124 ) , .B2( u0_u11_u6_n151 ) , .A2( u0_u11_u6_n93 ) );
  NAND4_X1 u0_u11_u6_U79 (.ZN( u0_out11_12 ) , .A4( u0_u11_u6_n114 ) , .A3( u0_u11_u6_n115 ) , .A2( u0_u11_u6_n116 ) , .A1( u0_u11_u6_n117 ) );
  AOI21_X1 u0_u11_u6_U8 (.B1( u0_u11_u6_n107 ) , .B2( u0_u11_u6_n132 ) , .A( u0_u11_u6_n158 ) , .ZN( u0_u11_u6_n88 ) );
  OAI22_X1 u0_u11_u6_U80 (.B2( u0_u11_u6_n111 ) , .ZN( u0_u11_u6_n116 ) , .B1( u0_u11_u6_n126 ) , .A2( u0_u11_u6_n164 ) , .A1( u0_u11_u6_n167 ) );
  OAI21_X1 u0_u11_u6_U81 (.A( u0_u11_u6_n108 ) , .ZN( u0_u11_u6_n117 ) , .B2( u0_u11_u6_n141 ) , .B1( u0_u11_u6_n163 ) );
  OAI211_X1 u0_u11_u6_U82 (.ZN( u0_out11_7 ) , .B( u0_u11_u6_n153 ) , .C2( u0_u11_u6_n154 ) , .C1( u0_u11_u6_n155 ) , .A( u0_u11_u6_n174 ) );
  NOR3_X1 u0_u11_u6_U83 (.A1( u0_u11_u6_n141 ) , .ZN( u0_u11_u6_n154 ) , .A3( u0_u11_u6_n164 ) , .A2( u0_u11_u6_n171 ) );
  AOI211_X1 u0_u11_u6_U84 (.B( u0_u11_u6_n149 ) , .A( u0_u11_u6_n150 ) , .C2( u0_u11_u6_n151 ) , .C1( u0_u11_u6_n152 ) , .ZN( u0_u11_u6_n153 ) );
  OAI211_X1 u0_u11_u6_U85 (.ZN( u0_out11_22 ) , .B( u0_u11_u6_n137 ) , .A( u0_u11_u6_n138 ) , .C2( u0_u11_u6_n139 ) , .C1( u0_u11_u6_n140 ) );
  AOI22_X1 u0_u11_u6_U86 (.B1( u0_u11_u6_n124 ) , .A2( u0_u11_u6_n125 ) , .A1( u0_u11_u6_n126 ) , .ZN( u0_u11_u6_n138 ) , .B2( u0_u11_u6_n161 ) );
  AND4_X1 u0_u11_u6_U87 (.A3( u0_u11_u6_n119 ) , .A1( u0_u11_u6_n120 ) , .A4( u0_u11_u6_n129 ) , .ZN( u0_u11_u6_n140 ) , .A2( u0_u11_u6_n143 ) );
  NAND3_X1 u0_u11_u6_U88 (.A2( u0_u11_u6_n123 ) , .ZN( u0_u11_u6_n125 ) , .A1( u0_u11_u6_n130 ) , .A3( u0_u11_u6_n131 ) );
  NAND3_X1 u0_u11_u6_U89 (.A3( u0_u11_u6_n133 ) , .ZN( u0_u11_u6_n141 ) , .A1( u0_u11_u6_n145 ) , .A2( u0_u11_u6_n148 ) );
  AOI21_X1 u0_u11_u6_U9 (.B2( u0_u11_u6_n147 ) , .B1( u0_u11_u6_n148 ) , .ZN( u0_u11_u6_n149 ) , .A( u0_u11_u6_n158 ) );
  NAND3_X1 u0_u11_u6_U90 (.ZN( u0_u11_u6_n101 ) , .A3( u0_u11_u6_n107 ) , .A2( u0_u11_u6_n121 ) , .A1( u0_u11_u6_n127 ) );
  NAND3_X1 u0_u11_u6_U91 (.ZN( u0_u11_u6_n102 ) , .A3( u0_u11_u6_n130 ) , .A2( u0_u11_u6_n145 ) , .A1( u0_u11_u6_n166 ) );
  NAND3_X1 u0_u11_u6_U92 (.A3( u0_u11_u6_n113 ) , .A1( u0_u11_u6_n119 ) , .A2( u0_u11_u6_n123 ) , .ZN( u0_u11_u6_n93 ) );
  NAND3_X1 u0_u11_u6_U93 (.ZN( u0_u11_u6_n142 ) , .A2( u0_u11_u6_n172 ) , .A3( u0_u11_u6_n89 ) , .A1( u0_u11_u6_n90 ) );
  AND3_X1 u0_u11_u7_U10 (.A3( u0_u11_u7_n110 ) , .A2( u0_u11_u7_n127 ) , .A1( u0_u11_u7_n132 ) , .ZN( u0_u11_u7_n92 ) );
  OAI21_X1 u0_u11_u7_U11 (.A( u0_u11_u7_n161 ) , .B1( u0_u11_u7_n168 ) , .B2( u0_u11_u7_n173 ) , .ZN( u0_u11_u7_n91 ) );
  AOI211_X1 u0_u11_u7_U12 (.A( u0_u11_u7_n117 ) , .ZN( u0_u11_u7_n118 ) , .C2( u0_u11_u7_n126 ) , .C1( u0_u11_u7_n177 ) , .B( u0_u11_u7_n180 ) );
  OAI22_X1 u0_u11_u7_U13 (.B1( u0_u11_u7_n115 ) , .ZN( u0_u11_u7_n117 ) , .A2( u0_u11_u7_n133 ) , .A1( u0_u11_u7_n137 ) , .B2( u0_u11_u7_n162 ) );
  INV_X1 u0_u11_u7_U14 (.A( u0_u11_u7_n116 ) , .ZN( u0_u11_u7_n180 ) );
  NOR3_X1 u0_u11_u7_U15 (.ZN( u0_u11_u7_n115 ) , .A3( u0_u11_u7_n145 ) , .A2( u0_u11_u7_n168 ) , .A1( u0_u11_u7_n169 ) );
  OAI211_X1 u0_u11_u7_U16 (.B( u0_u11_u7_n122 ) , .A( u0_u11_u7_n123 ) , .C2( u0_u11_u7_n124 ) , .ZN( u0_u11_u7_n154 ) , .C1( u0_u11_u7_n162 ) );
  AOI222_X1 u0_u11_u7_U17 (.ZN( u0_u11_u7_n122 ) , .C2( u0_u11_u7_n126 ) , .C1( u0_u11_u7_n145 ) , .B1( u0_u11_u7_n161 ) , .A2( u0_u11_u7_n165 ) , .B2( u0_u11_u7_n170 ) , .A1( u0_u11_u7_n176 ) );
  INV_X1 u0_u11_u7_U18 (.A( u0_u11_u7_n133 ) , .ZN( u0_u11_u7_n176 ) );
  NOR3_X1 u0_u11_u7_U19 (.A2( u0_u11_u7_n134 ) , .A1( u0_u11_u7_n135 ) , .ZN( u0_u11_u7_n136 ) , .A3( u0_u11_u7_n171 ) );
  NOR2_X1 u0_u11_u7_U20 (.A1( u0_u11_u7_n130 ) , .A2( u0_u11_u7_n134 ) , .ZN( u0_u11_u7_n153 ) );
  INV_X1 u0_u11_u7_U21 (.A( u0_u11_u7_n101 ) , .ZN( u0_u11_u7_n165 ) );
  NOR2_X1 u0_u11_u7_U22 (.ZN( u0_u11_u7_n111 ) , .A2( u0_u11_u7_n134 ) , .A1( u0_u11_u7_n169 ) );
  AOI21_X1 u0_u11_u7_U23 (.ZN( u0_u11_u7_n104 ) , .B2( u0_u11_u7_n112 ) , .B1( u0_u11_u7_n127 ) , .A( u0_u11_u7_n164 ) );
  AOI21_X1 u0_u11_u7_U24 (.ZN( u0_u11_u7_n106 ) , .B1( u0_u11_u7_n133 ) , .B2( u0_u11_u7_n146 ) , .A( u0_u11_u7_n162 ) );
  AOI21_X1 u0_u11_u7_U25 (.A( u0_u11_u7_n101 ) , .ZN( u0_u11_u7_n107 ) , .B2( u0_u11_u7_n128 ) , .B1( u0_u11_u7_n175 ) );
  INV_X1 u0_u11_u7_U26 (.A( u0_u11_u7_n138 ) , .ZN( u0_u11_u7_n171 ) );
  INV_X1 u0_u11_u7_U27 (.A( u0_u11_u7_n131 ) , .ZN( u0_u11_u7_n177 ) );
  INV_X1 u0_u11_u7_U28 (.A( u0_u11_u7_n110 ) , .ZN( u0_u11_u7_n174 ) );
  NAND2_X1 u0_u11_u7_U29 (.A1( u0_u11_u7_n129 ) , .A2( u0_u11_u7_n132 ) , .ZN( u0_u11_u7_n149 ) );
  OAI21_X1 u0_u11_u7_U3 (.ZN( u0_u11_u7_n159 ) , .A( u0_u11_u7_n165 ) , .B2( u0_u11_u7_n171 ) , .B1( u0_u11_u7_n174 ) );
  NAND2_X1 u0_u11_u7_U30 (.A1( u0_u11_u7_n113 ) , .A2( u0_u11_u7_n124 ) , .ZN( u0_u11_u7_n130 ) );
  INV_X1 u0_u11_u7_U31 (.A( u0_u11_u7_n112 ) , .ZN( u0_u11_u7_n173 ) );
  INV_X1 u0_u11_u7_U32 (.A( u0_u11_u7_n128 ) , .ZN( u0_u11_u7_n168 ) );
  INV_X1 u0_u11_u7_U33 (.A( u0_u11_u7_n148 ) , .ZN( u0_u11_u7_n169 ) );
  INV_X1 u0_u11_u7_U34 (.A( u0_u11_u7_n127 ) , .ZN( u0_u11_u7_n179 ) );
  NOR2_X1 u0_u11_u7_U35 (.ZN( u0_u11_u7_n101 ) , .A2( u0_u11_u7_n150 ) , .A1( u0_u11_u7_n156 ) );
  AOI211_X1 u0_u11_u7_U36 (.B( u0_u11_u7_n154 ) , .A( u0_u11_u7_n155 ) , .C1( u0_u11_u7_n156 ) , .ZN( u0_u11_u7_n157 ) , .C2( u0_u11_u7_n172 ) );
  INV_X1 u0_u11_u7_U37 (.A( u0_u11_u7_n153 ) , .ZN( u0_u11_u7_n172 ) );
  AOI211_X1 u0_u11_u7_U38 (.B( u0_u11_u7_n139 ) , .A( u0_u11_u7_n140 ) , .C2( u0_u11_u7_n141 ) , .ZN( u0_u11_u7_n142 ) , .C1( u0_u11_u7_n156 ) );
  AOI21_X1 u0_u11_u7_U39 (.A( u0_u11_u7_n137 ) , .B1( u0_u11_u7_n138 ) , .ZN( u0_u11_u7_n139 ) , .B2( u0_u11_u7_n146 ) );
  INV_X1 u0_u11_u7_U4 (.A( u0_u11_u7_n111 ) , .ZN( u0_u11_u7_n170 ) );
  NAND4_X1 u0_u11_u7_U40 (.A3( u0_u11_u7_n127 ) , .A2( u0_u11_u7_n128 ) , .A1( u0_u11_u7_n129 ) , .ZN( u0_u11_u7_n141 ) , .A4( u0_u11_u7_n147 ) );
  OAI22_X1 u0_u11_u7_U41 (.B1( u0_u11_u7_n136 ) , .ZN( u0_u11_u7_n140 ) , .A1( u0_u11_u7_n153 ) , .B2( u0_u11_u7_n162 ) , .A2( u0_u11_u7_n164 ) );
  AOI21_X1 u0_u11_u7_U42 (.ZN( u0_u11_u7_n123 ) , .B1( u0_u11_u7_n165 ) , .B2( u0_u11_u7_n177 ) , .A( u0_u11_u7_n97 ) );
  AOI21_X1 u0_u11_u7_U43 (.B2( u0_u11_u7_n113 ) , .B1( u0_u11_u7_n124 ) , .A( u0_u11_u7_n125 ) , .ZN( u0_u11_u7_n97 ) );
  INV_X1 u0_u11_u7_U44 (.A( u0_u11_u7_n125 ) , .ZN( u0_u11_u7_n161 ) );
  INV_X1 u0_u11_u7_U45 (.A( u0_u11_u7_n152 ) , .ZN( u0_u11_u7_n162 ) );
  AOI22_X1 u0_u11_u7_U46 (.A2( u0_u11_u7_n114 ) , .ZN( u0_u11_u7_n119 ) , .B1( u0_u11_u7_n130 ) , .A1( u0_u11_u7_n156 ) , .B2( u0_u11_u7_n165 ) );
  NAND2_X1 u0_u11_u7_U47 (.A2( u0_u11_u7_n112 ) , .ZN( u0_u11_u7_n114 ) , .A1( u0_u11_u7_n175 ) );
  AND2_X1 u0_u11_u7_U48 (.ZN( u0_u11_u7_n145 ) , .A2( u0_u11_u7_n98 ) , .A1( u0_u11_u7_n99 ) );
  NOR2_X1 u0_u11_u7_U49 (.ZN( u0_u11_u7_n137 ) , .A1( u0_u11_u7_n150 ) , .A2( u0_u11_u7_n161 ) );
  INV_X1 u0_u11_u7_U5 (.A( u0_u11_u7_n149 ) , .ZN( u0_u11_u7_n175 ) );
  AOI21_X1 u0_u11_u7_U50 (.ZN( u0_u11_u7_n105 ) , .B2( u0_u11_u7_n110 ) , .A( u0_u11_u7_n125 ) , .B1( u0_u11_u7_n147 ) );
  NAND2_X1 u0_u11_u7_U51 (.ZN( u0_u11_u7_n146 ) , .A1( u0_u11_u7_n95 ) , .A2( u0_u11_u7_n98 ) );
  NAND2_X1 u0_u11_u7_U52 (.A2( u0_u11_u7_n103 ) , .ZN( u0_u11_u7_n147 ) , .A1( u0_u11_u7_n93 ) );
  NAND2_X1 u0_u11_u7_U53 (.A1( u0_u11_u7_n103 ) , .ZN( u0_u11_u7_n127 ) , .A2( u0_u11_u7_n99 ) );
  OR2_X1 u0_u11_u7_U54 (.ZN( u0_u11_u7_n126 ) , .A2( u0_u11_u7_n152 ) , .A1( u0_u11_u7_n156 ) );
  NAND2_X1 u0_u11_u7_U55 (.A2( u0_u11_u7_n102 ) , .A1( u0_u11_u7_n103 ) , .ZN( u0_u11_u7_n133 ) );
  NAND2_X1 u0_u11_u7_U56 (.ZN( u0_u11_u7_n112 ) , .A2( u0_u11_u7_n96 ) , .A1( u0_u11_u7_n99 ) );
  NAND2_X1 u0_u11_u7_U57 (.A2( u0_u11_u7_n102 ) , .ZN( u0_u11_u7_n128 ) , .A1( u0_u11_u7_n98 ) );
  NAND2_X1 u0_u11_u7_U58 (.A1( u0_u11_u7_n100 ) , .ZN( u0_u11_u7_n113 ) , .A2( u0_u11_u7_n93 ) );
  NAND2_X1 u0_u11_u7_U59 (.A2( u0_u11_u7_n102 ) , .ZN( u0_u11_u7_n124 ) , .A1( u0_u11_u7_n96 ) );
  INV_X1 u0_u11_u7_U6 (.A( u0_u11_u7_n154 ) , .ZN( u0_u11_u7_n178 ) );
  NAND2_X1 u0_u11_u7_U60 (.ZN( u0_u11_u7_n110 ) , .A1( u0_u11_u7_n95 ) , .A2( u0_u11_u7_n96 ) );
  INV_X1 u0_u11_u7_U61 (.A( u0_u11_u7_n150 ) , .ZN( u0_u11_u7_n164 ) );
  AND2_X1 u0_u11_u7_U62 (.ZN( u0_u11_u7_n134 ) , .A1( u0_u11_u7_n93 ) , .A2( u0_u11_u7_n98 ) );
  NAND2_X1 u0_u11_u7_U63 (.A1( u0_u11_u7_n100 ) , .A2( u0_u11_u7_n102 ) , .ZN( u0_u11_u7_n129 ) );
  NAND2_X1 u0_u11_u7_U64 (.A2( u0_u11_u7_n103 ) , .ZN( u0_u11_u7_n131 ) , .A1( u0_u11_u7_n95 ) );
  NAND2_X1 u0_u11_u7_U65 (.A1( u0_u11_u7_n100 ) , .ZN( u0_u11_u7_n138 ) , .A2( u0_u11_u7_n99 ) );
  NAND2_X1 u0_u11_u7_U66 (.ZN( u0_u11_u7_n132 ) , .A1( u0_u11_u7_n93 ) , .A2( u0_u11_u7_n96 ) );
  NAND2_X1 u0_u11_u7_U67 (.A1( u0_u11_u7_n100 ) , .ZN( u0_u11_u7_n148 ) , .A2( u0_u11_u7_n95 ) );
  NOR2_X1 u0_u11_u7_U68 (.A2( u0_u11_X_47 ) , .ZN( u0_u11_u7_n150 ) , .A1( u0_u11_u7_n163 ) );
  NOR2_X1 u0_u11_u7_U69 (.A2( u0_u11_X_43 ) , .A1( u0_u11_X_44 ) , .ZN( u0_u11_u7_n103 ) );
  AOI211_X1 u0_u11_u7_U7 (.ZN( u0_u11_u7_n116 ) , .A( u0_u11_u7_n155 ) , .C1( u0_u11_u7_n161 ) , .C2( u0_u11_u7_n171 ) , .B( u0_u11_u7_n94 ) );
  NOR2_X1 u0_u11_u7_U70 (.A2( u0_u11_X_48 ) , .A1( u0_u11_u7_n166 ) , .ZN( u0_u11_u7_n95 ) );
  NOR2_X1 u0_u11_u7_U71 (.A2( u0_u11_X_45 ) , .A1( u0_u11_X_48 ) , .ZN( u0_u11_u7_n99 ) );
  NOR2_X1 u0_u11_u7_U72 (.A2( u0_u11_X_44 ) , .A1( u0_u11_u7_n167 ) , .ZN( u0_u11_u7_n98 ) );
  NOR2_X1 u0_u11_u7_U73 (.A2( u0_u11_X_46 ) , .A1( u0_u11_X_47 ) , .ZN( u0_u11_u7_n152 ) );
  AND2_X1 u0_u11_u7_U74 (.A1( u0_u11_X_47 ) , .ZN( u0_u11_u7_n156 ) , .A2( u0_u11_u7_n163 ) );
  NAND2_X1 u0_u11_u7_U75 (.A2( u0_u11_X_46 ) , .A1( u0_u11_X_47 ) , .ZN( u0_u11_u7_n125 ) );
  AND2_X1 u0_u11_u7_U76 (.A2( u0_u11_X_45 ) , .A1( u0_u11_X_48 ) , .ZN( u0_u11_u7_n102 ) );
  AND2_X1 u0_u11_u7_U77 (.A2( u0_u11_X_43 ) , .A1( u0_u11_X_44 ) , .ZN( u0_u11_u7_n96 ) );
  AND2_X1 u0_u11_u7_U78 (.A1( u0_u11_X_44 ) , .ZN( u0_u11_u7_n100 ) , .A2( u0_u11_u7_n167 ) );
  AND2_X1 u0_u11_u7_U79 (.A1( u0_u11_X_48 ) , .A2( u0_u11_u7_n166 ) , .ZN( u0_u11_u7_n93 ) );
  OAI222_X1 u0_u11_u7_U8 (.C2( u0_u11_u7_n101 ) , .B2( u0_u11_u7_n111 ) , .A1( u0_u11_u7_n113 ) , .C1( u0_u11_u7_n146 ) , .A2( u0_u11_u7_n162 ) , .B1( u0_u11_u7_n164 ) , .ZN( u0_u11_u7_n94 ) );
  INV_X1 u0_u11_u7_U80 (.A( u0_u11_X_46 ) , .ZN( u0_u11_u7_n163 ) );
  INV_X1 u0_u11_u7_U81 (.A( u0_u11_X_43 ) , .ZN( u0_u11_u7_n167 ) );
  INV_X1 u0_u11_u7_U82 (.A( u0_u11_X_45 ) , .ZN( u0_u11_u7_n166 ) );
  NAND4_X1 u0_u11_u7_U83 (.ZN( u0_out11_27 ) , .A4( u0_u11_u7_n118 ) , .A3( u0_u11_u7_n119 ) , .A2( u0_u11_u7_n120 ) , .A1( u0_u11_u7_n121 ) );
  OAI21_X1 u0_u11_u7_U84 (.ZN( u0_u11_u7_n121 ) , .B2( u0_u11_u7_n145 ) , .A( u0_u11_u7_n150 ) , .B1( u0_u11_u7_n174 ) );
  OAI21_X1 u0_u11_u7_U85 (.ZN( u0_u11_u7_n120 ) , .A( u0_u11_u7_n161 ) , .B2( u0_u11_u7_n170 ) , .B1( u0_u11_u7_n179 ) );
  NAND4_X1 u0_u11_u7_U86 (.ZN( u0_out11_21 ) , .A4( u0_u11_u7_n157 ) , .A3( u0_u11_u7_n158 ) , .A2( u0_u11_u7_n159 ) , .A1( u0_u11_u7_n160 ) );
  OAI21_X1 u0_u11_u7_U87 (.B1( u0_u11_u7_n145 ) , .ZN( u0_u11_u7_n160 ) , .A( u0_u11_u7_n161 ) , .B2( u0_u11_u7_n177 ) );
  AOI22_X1 u0_u11_u7_U88 (.B2( u0_u11_u7_n149 ) , .B1( u0_u11_u7_n150 ) , .A2( u0_u11_u7_n151 ) , .A1( u0_u11_u7_n152 ) , .ZN( u0_u11_u7_n158 ) );
  NAND4_X1 u0_u11_u7_U89 (.ZN( u0_out11_15 ) , .A4( u0_u11_u7_n142 ) , .A3( u0_u11_u7_n143 ) , .A2( u0_u11_u7_n144 ) , .A1( u0_u11_u7_n178 ) );
  OAI221_X1 u0_u11_u7_U9 (.C1( u0_u11_u7_n101 ) , .C2( u0_u11_u7_n147 ) , .ZN( u0_u11_u7_n155 ) , .B2( u0_u11_u7_n162 ) , .A( u0_u11_u7_n91 ) , .B1( u0_u11_u7_n92 ) );
  OR2_X1 u0_u11_u7_U90 (.A2( u0_u11_u7_n125 ) , .A1( u0_u11_u7_n129 ) , .ZN( u0_u11_u7_n144 ) );
  AOI22_X1 u0_u11_u7_U91 (.A2( u0_u11_u7_n126 ) , .ZN( u0_u11_u7_n143 ) , .B2( u0_u11_u7_n165 ) , .B1( u0_u11_u7_n173 ) , .A1( u0_u11_u7_n174 ) );
  NAND4_X1 u0_u11_u7_U92 (.ZN( u0_out11_5 ) , .A4( u0_u11_u7_n108 ) , .A3( u0_u11_u7_n109 ) , .A1( u0_u11_u7_n116 ) , .A2( u0_u11_u7_n123 ) );
  AOI22_X1 u0_u11_u7_U93 (.ZN( u0_u11_u7_n109 ) , .A2( u0_u11_u7_n126 ) , .B2( u0_u11_u7_n145 ) , .B1( u0_u11_u7_n156 ) , .A1( u0_u11_u7_n171 ) );
  NOR4_X1 u0_u11_u7_U94 (.A4( u0_u11_u7_n104 ) , .A3( u0_u11_u7_n105 ) , .A2( u0_u11_u7_n106 ) , .A1( u0_u11_u7_n107 ) , .ZN( u0_u11_u7_n108 ) );
  NAND3_X1 u0_u11_u7_U95 (.A3( u0_u11_u7_n146 ) , .A2( u0_u11_u7_n147 ) , .A1( u0_u11_u7_n148 ) , .ZN( u0_u11_u7_n151 ) );
  NAND3_X1 u0_u11_u7_U96 (.A3( u0_u11_u7_n131 ) , .A2( u0_u11_u7_n132 ) , .A1( u0_u11_u7_n133 ) , .ZN( u0_u11_u7_n135 ) );
  XOR2_X1 u0_u12_U10 (.B( u0_K13_45 ) , .A( u0_R11_30 ) , .Z( u0_u12_X_45 ) );
  XOR2_X1 u0_u12_U11 (.B( u0_K13_44 ) , .A( u0_R11_29 ) , .Z( u0_u12_X_44 ) );
  XOR2_X1 u0_u12_U12 (.B( u0_K13_43 ) , .A( u0_R11_28 ) , .Z( u0_u12_X_43 ) );
  XOR2_X1 u0_u12_U16 (.B( u0_K13_3 ) , .A( u0_R11_2 ) , .Z( u0_u12_X_3 ) );
  XOR2_X1 u0_u12_U27 (.B( u0_K13_2 ) , .A( u0_R11_1 ) , .Z( u0_u12_X_2 ) );
  XOR2_X1 u0_u12_U38 (.B( u0_K13_1 ) , .A( u0_R11_32 ) , .Z( u0_u12_X_1 ) );
  XOR2_X1 u0_u12_U4 (.B( u0_K13_6 ) , .A( u0_R11_5 ) , .Z( u0_u12_X_6 ) );
  XOR2_X1 u0_u12_U5 (.B( u0_K13_5 ) , .A( u0_R11_4 ) , .Z( u0_u12_X_5 ) );
  XOR2_X1 u0_u12_U6 (.B( u0_K13_4 ) , .A( u0_R11_3 ) , .Z( u0_u12_X_4 ) );
  XOR2_X1 u0_u12_U7 (.B( u0_K13_48 ) , .A( u0_R11_1 ) , .Z( u0_u12_X_48 ) );
  XOR2_X1 u0_u12_U8 (.B( u0_K13_47 ) , .A( u0_R11_32 ) , .Z( u0_u12_X_47 ) );
  XOR2_X1 u0_u12_U9 (.B( u0_K13_46 ) , .A( u0_R11_31 ) , .Z( u0_u12_X_46 ) );
  NAND2_X1 u0_u12_u0_U10 (.ZN( u0_u12_u0_n113 ) , .A1( u0_u12_u0_n139 ) , .A2( u0_u12_u0_n149 ) );
  AND3_X1 u0_u12_u0_U11 (.A2( u0_u12_u0_n112 ) , .ZN( u0_u12_u0_n127 ) , .A3( u0_u12_u0_n130 ) , .A1( u0_u12_u0_n148 ) );
  AND2_X1 u0_u12_u0_U12 (.ZN( u0_u12_u0_n107 ) , .A1( u0_u12_u0_n130 ) , .A2( u0_u12_u0_n140 ) );
  AND2_X1 u0_u12_u0_U13 (.A2( u0_u12_u0_n129 ) , .A1( u0_u12_u0_n130 ) , .ZN( u0_u12_u0_n151 ) );
  AND2_X1 u0_u12_u0_U14 (.A1( u0_u12_u0_n108 ) , .A2( u0_u12_u0_n125 ) , .ZN( u0_u12_u0_n145 ) );
  INV_X1 u0_u12_u0_U15 (.A( u0_u12_u0_n143 ) , .ZN( u0_u12_u0_n173 ) );
  NOR2_X1 u0_u12_u0_U16 (.A2( u0_u12_u0_n136 ) , .ZN( u0_u12_u0_n147 ) , .A1( u0_u12_u0_n160 ) );
  AOI21_X1 u0_u12_u0_U17 (.B1( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n132 ) , .A( u0_u12_u0_n165 ) , .B2( u0_u12_u0_n93 ) );
  INV_X1 u0_u12_u0_U18 (.A( u0_u12_u0_n142 ) , .ZN( u0_u12_u0_n165 ) );
  OAI22_X1 u0_u12_u0_U19 (.B1( u0_u12_u0_n131 ) , .A1( u0_u12_u0_n144 ) , .B2( u0_u12_u0_n147 ) , .A2( u0_u12_u0_n90 ) , .ZN( u0_u12_u0_n91 ) );
  AND3_X1 u0_u12_u0_U20 (.A3( u0_u12_u0_n121 ) , .A2( u0_u12_u0_n125 ) , .A1( u0_u12_u0_n148 ) , .ZN( u0_u12_u0_n90 ) );
  OAI22_X1 u0_u12_u0_U21 (.B1( u0_u12_u0_n125 ) , .ZN( u0_u12_u0_n126 ) , .A1( u0_u12_u0_n138 ) , .A2( u0_u12_u0_n146 ) , .B2( u0_u12_u0_n147 ) );
  INV_X1 u0_u12_u0_U22 (.A( u0_u12_u0_n136 ) , .ZN( u0_u12_u0_n161 ) );
  AOI22_X1 u0_u12_u0_U23 (.B2( u0_u12_u0_n109 ) , .A2( u0_u12_u0_n110 ) , .ZN( u0_u12_u0_n111 ) , .B1( u0_u12_u0_n118 ) , .A1( u0_u12_u0_n160 ) );
  NAND2_X1 u0_u12_u0_U24 (.A2( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n140 ) , .A1( u0_u12_u0_n94 ) );
  NAND2_X1 u0_u12_u0_U25 (.A2( u0_u12_u0_n102 ) , .A1( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n149 ) );
  INV_X1 u0_u12_u0_U26 (.A( u0_u12_u0_n118 ) , .ZN( u0_u12_u0_n158 ) );
  NAND2_X1 u0_u12_u0_U27 (.A2( u0_u12_u0_n100 ) , .ZN( u0_u12_u0_n131 ) , .A1( u0_u12_u0_n92 ) );
  NAND2_X1 u0_u12_u0_U28 (.ZN( u0_u12_u0_n108 ) , .A1( u0_u12_u0_n92 ) , .A2( u0_u12_u0_n94 ) );
  AOI21_X1 u0_u12_u0_U29 (.ZN( u0_u12_u0_n104 ) , .B1( u0_u12_u0_n107 ) , .B2( u0_u12_u0_n141 ) , .A( u0_u12_u0_n144 ) );
  INV_X1 u0_u12_u0_U3 (.A( u0_u12_u0_n113 ) , .ZN( u0_u12_u0_n166 ) );
  AOI21_X1 u0_u12_u0_U30 (.ZN( u0_u12_u0_n116 ) , .B2( u0_u12_u0_n142 ) , .A( u0_u12_u0_n144 ) , .B1( u0_u12_u0_n166 ) );
  AOI21_X1 u0_u12_u0_U31 (.B1( u0_u12_u0_n127 ) , .B2( u0_u12_u0_n129 ) , .A( u0_u12_u0_n138 ) , .ZN( u0_u12_u0_n96 ) );
  NAND2_X1 u0_u12_u0_U32 (.A2( u0_u12_u0_n102 ) , .ZN( u0_u12_u0_n114 ) , .A1( u0_u12_u0_n92 ) );
  NOR2_X1 u0_u12_u0_U33 (.A1( u0_u12_u0_n120 ) , .ZN( u0_u12_u0_n143 ) , .A2( u0_u12_u0_n167 ) );
  OAI221_X1 u0_u12_u0_U34 (.C1( u0_u12_u0_n112 ) , .ZN( u0_u12_u0_n120 ) , .B1( u0_u12_u0_n138 ) , .B2( u0_u12_u0_n141 ) , .C2( u0_u12_u0_n147 ) , .A( u0_u12_u0_n172 ) );
  AOI211_X1 u0_u12_u0_U35 (.B( u0_u12_u0_n115 ) , .A( u0_u12_u0_n116 ) , .C2( u0_u12_u0_n117 ) , .C1( u0_u12_u0_n118 ) , .ZN( u0_u12_u0_n119 ) );
  NAND2_X1 u0_u12_u0_U36 (.A1( u0_u12_u0_n100 ) , .A2( u0_u12_u0_n103 ) , .ZN( u0_u12_u0_n125 ) );
  NAND2_X1 u0_u12_u0_U37 (.A1( u0_u12_u0_n101 ) , .A2( u0_u12_u0_n102 ) , .ZN( u0_u12_u0_n150 ) );
  INV_X1 u0_u12_u0_U38 (.A( u0_u12_u0_n138 ) , .ZN( u0_u12_u0_n160 ) );
  NAND2_X1 u0_u12_u0_U39 (.A2( u0_u12_u0_n100 ) , .A1( u0_u12_u0_n101 ) , .ZN( u0_u12_u0_n139 ) );
  AOI21_X1 u0_u12_u0_U4 (.B1( u0_u12_u0_n114 ) , .ZN( u0_u12_u0_n115 ) , .B2( u0_u12_u0_n129 ) , .A( u0_u12_u0_n161 ) );
  NAND2_X1 u0_u12_u0_U40 (.A1( u0_u12_u0_n101 ) , .ZN( u0_u12_u0_n130 ) , .A2( u0_u12_u0_n94 ) );
  NAND2_X1 u0_u12_u0_U41 (.ZN( u0_u12_u0_n112 ) , .A2( u0_u12_u0_n92 ) , .A1( u0_u12_u0_n93 ) );
  INV_X1 u0_u12_u0_U42 (.ZN( u0_u12_u0_n172 ) , .A( u0_u12_u0_n88 ) );
  OAI222_X1 u0_u12_u0_U43 (.C1( u0_u12_u0_n108 ) , .A1( u0_u12_u0_n125 ) , .B2( u0_u12_u0_n128 ) , .B1( u0_u12_u0_n144 ) , .A2( u0_u12_u0_n158 ) , .C2( u0_u12_u0_n161 ) , .ZN( u0_u12_u0_n88 ) );
  NAND2_X1 u0_u12_u0_U44 (.A2( u0_u12_u0_n101 ) , .ZN( u0_u12_u0_n121 ) , .A1( u0_u12_u0_n93 ) );
  OR3_X1 u0_u12_u0_U45 (.A3( u0_u12_u0_n152 ) , .A2( u0_u12_u0_n153 ) , .A1( u0_u12_u0_n154 ) , .ZN( u0_u12_u0_n155 ) );
  AOI21_X1 u0_u12_u0_U46 (.A( u0_u12_u0_n144 ) , .B2( u0_u12_u0_n145 ) , .B1( u0_u12_u0_n146 ) , .ZN( u0_u12_u0_n154 ) );
  AOI21_X1 u0_u12_u0_U47 (.B2( u0_u12_u0_n150 ) , .B1( u0_u12_u0_n151 ) , .ZN( u0_u12_u0_n152 ) , .A( u0_u12_u0_n158 ) );
  AOI21_X1 u0_u12_u0_U48 (.A( u0_u12_u0_n147 ) , .B2( u0_u12_u0_n148 ) , .B1( u0_u12_u0_n149 ) , .ZN( u0_u12_u0_n153 ) );
  INV_X1 u0_u12_u0_U49 (.ZN( u0_u12_u0_n171 ) , .A( u0_u12_u0_n99 ) );
  AOI21_X1 u0_u12_u0_U5 (.B2( u0_u12_u0_n131 ) , .ZN( u0_u12_u0_n134 ) , .B1( u0_u12_u0_n151 ) , .A( u0_u12_u0_n158 ) );
  OAI211_X1 u0_u12_u0_U50 (.C2( u0_u12_u0_n140 ) , .C1( u0_u12_u0_n161 ) , .A( u0_u12_u0_n169 ) , .B( u0_u12_u0_n98 ) , .ZN( u0_u12_u0_n99 ) );
  INV_X1 u0_u12_u0_U51 (.ZN( u0_u12_u0_n169 ) , .A( u0_u12_u0_n91 ) );
  AOI211_X1 u0_u12_u0_U52 (.C1( u0_u12_u0_n118 ) , .A( u0_u12_u0_n123 ) , .B( u0_u12_u0_n96 ) , .C2( u0_u12_u0_n97 ) , .ZN( u0_u12_u0_n98 ) );
  NOR2_X1 u0_u12_u0_U53 (.A2( u0_u12_X_4 ) , .A1( u0_u12_X_5 ) , .ZN( u0_u12_u0_n118 ) );
  NOR2_X1 u0_u12_u0_U54 (.A2( u0_u12_X_1 ) , .ZN( u0_u12_u0_n101 ) , .A1( u0_u12_u0_n163 ) );
  NOR2_X1 u0_u12_u0_U55 (.A2( u0_u12_X_6 ) , .ZN( u0_u12_u0_n100 ) , .A1( u0_u12_u0_n162 ) );
  NAND2_X1 u0_u12_u0_U56 (.A2( u0_u12_X_4 ) , .A1( u0_u12_X_5 ) , .ZN( u0_u12_u0_n144 ) );
  NOR2_X1 u0_u12_u0_U57 (.A2( u0_u12_X_5 ) , .ZN( u0_u12_u0_n136 ) , .A1( u0_u12_u0_n159 ) );
  NAND2_X1 u0_u12_u0_U58 (.A1( u0_u12_X_5 ) , .ZN( u0_u12_u0_n138 ) , .A2( u0_u12_u0_n159 ) );
  AND2_X1 u0_u12_u0_U59 (.A2( u0_u12_X_3 ) , .A1( u0_u12_X_6 ) , .ZN( u0_u12_u0_n102 ) );
  NOR2_X1 u0_u12_u0_U6 (.A1( u0_u12_u0_n108 ) , .ZN( u0_u12_u0_n123 ) , .A2( u0_u12_u0_n158 ) );
  AND2_X1 u0_u12_u0_U60 (.A1( u0_u12_X_6 ) , .A2( u0_u12_u0_n162 ) , .ZN( u0_u12_u0_n93 ) );
  INV_X1 u0_u12_u0_U61 (.A( u0_u12_X_4 ) , .ZN( u0_u12_u0_n159 ) );
  INV_X1 u0_u12_u0_U62 (.A( u0_u12_X_3 ) , .ZN( u0_u12_u0_n162 ) );
  INV_X1 u0_u12_u0_U63 (.A( u0_u12_u0_n126 ) , .ZN( u0_u12_u0_n168 ) );
  AOI211_X1 u0_u12_u0_U64 (.B( u0_u12_u0_n133 ) , .A( u0_u12_u0_n134 ) , .C2( u0_u12_u0_n135 ) , .C1( u0_u12_u0_n136 ) , .ZN( u0_u12_u0_n137 ) );
  OR4_X1 u0_u12_u0_U65 (.ZN( u0_out12_17 ) , .A4( u0_u12_u0_n122 ) , .A2( u0_u12_u0_n123 ) , .A1( u0_u12_u0_n124 ) , .A3( u0_u12_u0_n170 ) );
  AOI21_X1 u0_u12_u0_U66 (.B2( u0_u12_u0_n107 ) , .ZN( u0_u12_u0_n124 ) , .B1( u0_u12_u0_n128 ) , .A( u0_u12_u0_n161 ) );
  INV_X1 u0_u12_u0_U67 (.A( u0_u12_u0_n111 ) , .ZN( u0_u12_u0_n170 ) );
  OR4_X1 u0_u12_u0_U68 (.ZN( u0_out12_31 ) , .A4( u0_u12_u0_n155 ) , .A2( u0_u12_u0_n156 ) , .A1( u0_u12_u0_n157 ) , .A3( u0_u12_u0_n173 ) );
  AOI21_X1 u0_u12_u0_U69 (.A( u0_u12_u0_n138 ) , .B2( u0_u12_u0_n139 ) , .B1( u0_u12_u0_n140 ) , .ZN( u0_u12_u0_n157 ) );
  OAI21_X1 u0_u12_u0_U7 (.B1( u0_u12_u0_n150 ) , .B2( u0_u12_u0_n158 ) , .A( u0_u12_u0_n172 ) , .ZN( u0_u12_u0_n89 ) );
  AOI21_X1 u0_u12_u0_U70 (.B2( u0_u12_u0_n141 ) , .B1( u0_u12_u0_n142 ) , .ZN( u0_u12_u0_n156 ) , .A( u0_u12_u0_n161 ) );
  INV_X1 u0_u12_u0_U71 (.ZN( u0_u12_u0_n174 ) , .A( u0_u12_u0_n89 ) );
  AOI211_X1 u0_u12_u0_U72 (.B( u0_u12_u0_n104 ) , .A( u0_u12_u0_n105 ) , .ZN( u0_u12_u0_n106 ) , .C2( u0_u12_u0_n113 ) , .C1( u0_u12_u0_n160 ) );
  AND2_X1 u0_u12_u0_U73 (.A2( u0_u12_X_1 ) , .A1( u0_u12_X_2 ) , .ZN( u0_u12_u0_n95 ) );
  INV_X1 u0_u12_u0_U74 (.A( u0_u12_X_1 ) , .ZN( u0_u12_u0_n164 ) );
  NOR2_X1 u0_u12_u0_U75 (.A2( u0_u12_X_3 ) , .A1( u0_u12_X_6 ) , .ZN( u0_u12_u0_n94 ) );
  OAI221_X1 u0_u12_u0_U76 (.C1( u0_u12_u0_n121 ) , .ZN( u0_u12_u0_n122 ) , .B2( u0_u12_u0_n127 ) , .A( u0_u12_u0_n143 ) , .B1( u0_u12_u0_n144 ) , .C2( u0_u12_u0_n147 ) );
  AOI21_X1 u0_u12_u0_U77 (.B1( u0_u12_u0_n132 ) , .ZN( u0_u12_u0_n133 ) , .A( u0_u12_u0_n144 ) , .B2( u0_u12_u0_n166 ) );
  OAI22_X1 u0_u12_u0_U78 (.ZN( u0_u12_u0_n105 ) , .A2( u0_u12_u0_n132 ) , .B1( u0_u12_u0_n146 ) , .A1( u0_u12_u0_n147 ) , .B2( u0_u12_u0_n161 ) );
  NAND2_X1 u0_u12_u0_U79 (.ZN( u0_u12_u0_n110 ) , .A2( u0_u12_u0_n132 ) , .A1( u0_u12_u0_n145 ) );
  AND2_X1 u0_u12_u0_U8 (.A1( u0_u12_u0_n114 ) , .A2( u0_u12_u0_n121 ) , .ZN( u0_u12_u0_n146 ) );
  INV_X1 u0_u12_u0_U80 (.A( u0_u12_u0_n119 ) , .ZN( u0_u12_u0_n167 ) );
  NAND2_X1 u0_u12_u0_U81 (.ZN( u0_u12_u0_n148 ) , .A1( u0_u12_u0_n93 ) , .A2( u0_u12_u0_n95 ) );
  NAND2_X1 u0_u12_u0_U82 (.A1( u0_u12_u0_n100 ) , .ZN( u0_u12_u0_n129 ) , .A2( u0_u12_u0_n95 ) );
  NAND2_X1 u0_u12_u0_U83 (.A1( u0_u12_u0_n102 ) , .ZN( u0_u12_u0_n128 ) , .A2( u0_u12_u0_n95 ) );
  NOR2_X1 u0_u12_u0_U84 (.A2( u0_u12_X_1 ) , .A1( u0_u12_X_2 ) , .ZN( u0_u12_u0_n92 ) );
  NAND2_X1 u0_u12_u0_U85 (.ZN( u0_u12_u0_n142 ) , .A1( u0_u12_u0_n94 ) , .A2( u0_u12_u0_n95 ) );
  NOR2_X1 u0_u12_u0_U86 (.A2( u0_u12_X_2 ) , .ZN( u0_u12_u0_n103 ) , .A1( u0_u12_u0_n164 ) );
  INV_X1 u0_u12_u0_U87 (.A( u0_u12_X_2 ) , .ZN( u0_u12_u0_n163 ) );
  NAND3_X1 u0_u12_u0_U88 (.ZN( u0_out12_23 ) , .A3( u0_u12_u0_n137 ) , .A1( u0_u12_u0_n168 ) , .A2( u0_u12_u0_n171 ) );
  NAND3_X1 u0_u12_u0_U89 (.A3( u0_u12_u0_n127 ) , .A2( u0_u12_u0_n128 ) , .ZN( u0_u12_u0_n135 ) , .A1( u0_u12_u0_n150 ) );
  AND2_X1 u0_u12_u0_U9 (.A1( u0_u12_u0_n131 ) , .ZN( u0_u12_u0_n141 ) , .A2( u0_u12_u0_n150 ) );
  NAND3_X1 u0_u12_u0_U90 (.ZN( u0_u12_u0_n117 ) , .A3( u0_u12_u0_n132 ) , .A2( u0_u12_u0_n139 ) , .A1( u0_u12_u0_n148 ) );
  NAND3_X1 u0_u12_u0_U91 (.ZN( u0_u12_u0_n109 ) , .A2( u0_u12_u0_n114 ) , .A3( u0_u12_u0_n140 ) , .A1( u0_u12_u0_n149 ) );
  NAND3_X1 u0_u12_u0_U92 (.ZN( u0_out12_9 ) , .A3( u0_u12_u0_n106 ) , .A2( u0_u12_u0_n171 ) , .A1( u0_u12_u0_n174 ) );
  NAND3_X1 u0_u12_u0_U93 (.A2( u0_u12_u0_n128 ) , .A1( u0_u12_u0_n132 ) , .A3( u0_u12_u0_n146 ) , .ZN( u0_u12_u0_n97 ) );
  AND3_X1 u0_u12_u7_U10 (.A3( u0_u12_u7_n110 ) , .A2( u0_u12_u7_n127 ) , .A1( u0_u12_u7_n132 ) , .ZN( u0_u12_u7_n92 ) );
  OAI21_X1 u0_u12_u7_U11 (.A( u0_u12_u7_n161 ) , .B1( u0_u12_u7_n168 ) , .B2( u0_u12_u7_n173 ) , .ZN( u0_u12_u7_n91 ) );
  AOI211_X1 u0_u12_u7_U12 (.A( u0_u12_u7_n117 ) , .ZN( u0_u12_u7_n118 ) , .C2( u0_u12_u7_n126 ) , .C1( u0_u12_u7_n177 ) , .B( u0_u12_u7_n180 ) );
  OAI22_X1 u0_u12_u7_U13 (.B1( u0_u12_u7_n115 ) , .ZN( u0_u12_u7_n117 ) , .A2( u0_u12_u7_n133 ) , .A1( u0_u12_u7_n137 ) , .B2( u0_u12_u7_n162 ) );
  INV_X1 u0_u12_u7_U14 (.A( u0_u12_u7_n116 ) , .ZN( u0_u12_u7_n180 ) );
  NOR3_X1 u0_u12_u7_U15 (.ZN( u0_u12_u7_n115 ) , .A3( u0_u12_u7_n145 ) , .A2( u0_u12_u7_n168 ) , .A1( u0_u12_u7_n169 ) );
  OAI211_X1 u0_u12_u7_U16 (.B( u0_u12_u7_n122 ) , .A( u0_u12_u7_n123 ) , .C2( u0_u12_u7_n124 ) , .ZN( u0_u12_u7_n154 ) , .C1( u0_u12_u7_n162 ) );
  AOI222_X1 u0_u12_u7_U17 (.ZN( u0_u12_u7_n122 ) , .C2( u0_u12_u7_n126 ) , .C1( u0_u12_u7_n145 ) , .B1( u0_u12_u7_n161 ) , .A2( u0_u12_u7_n165 ) , .B2( u0_u12_u7_n170 ) , .A1( u0_u12_u7_n176 ) );
  INV_X1 u0_u12_u7_U18 (.A( u0_u12_u7_n133 ) , .ZN( u0_u12_u7_n176 ) );
  NOR3_X1 u0_u12_u7_U19 (.A2( u0_u12_u7_n134 ) , .A1( u0_u12_u7_n135 ) , .ZN( u0_u12_u7_n136 ) , .A3( u0_u12_u7_n171 ) );
  NOR2_X1 u0_u12_u7_U20 (.A1( u0_u12_u7_n130 ) , .A2( u0_u12_u7_n134 ) , .ZN( u0_u12_u7_n153 ) );
  INV_X1 u0_u12_u7_U21 (.A( u0_u12_u7_n101 ) , .ZN( u0_u12_u7_n165 ) );
  NOR2_X1 u0_u12_u7_U22 (.ZN( u0_u12_u7_n111 ) , .A2( u0_u12_u7_n134 ) , .A1( u0_u12_u7_n169 ) );
  AOI21_X1 u0_u12_u7_U23 (.ZN( u0_u12_u7_n104 ) , .B2( u0_u12_u7_n112 ) , .B1( u0_u12_u7_n127 ) , .A( u0_u12_u7_n164 ) );
  AOI21_X1 u0_u12_u7_U24 (.ZN( u0_u12_u7_n106 ) , .B1( u0_u12_u7_n133 ) , .B2( u0_u12_u7_n146 ) , .A( u0_u12_u7_n162 ) );
  AOI21_X1 u0_u12_u7_U25 (.A( u0_u12_u7_n101 ) , .ZN( u0_u12_u7_n107 ) , .B2( u0_u12_u7_n128 ) , .B1( u0_u12_u7_n175 ) );
  INV_X1 u0_u12_u7_U26 (.A( u0_u12_u7_n138 ) , .ZN( u0_u12_u7_n171 ) );
  INV_X1 u0_u12_u7_U27 (.A( u0_u12_u7_n131 ) , .ZN( u0_u12_u7_n177 ) );
  INV_X1 u0_u12_u7_U28 (.A( u0_u12_u7_n110 ) , .ZN( u0_u12_u7_n174 ) );
  NAND2_X1 u0_u12_u7_U29 (.A1( u0_u12_u7_n129 ) , .A2( u0_u12_u7_n132 ) , .ZN( u0_u12_u7_n149 ) );
  OAI21_X1 u0_u12_u7_U3 (.ZN( u0_u12_u7_n159 ) , .A( u0_u12_u7_n165 ) , .B2( u0_u12_u7_n171 ) , .B1( u0_u12_u7_n174 ) );
  NAND2_X1 u0_u12_u7_U30 (.A1( u0_u12_u7_n113 ) , .A2( u0_u12_u7_n124 ) , .ZN( u0_u12_u7_n130 ) );
  INV_X1 u0_u12_u7_U31 (.A( u0_u12_u7_n112 ) , .ZN( u0_u12_u7_n173 ) );
  INV_X1 u0_u12_u7_U32 (.A( u0_u12_u7_n128 ) , .ZN( u0_u12_u7_n168 ) );
  INV_X1 u0_u12_u7_U33 (.A( u0_u12_u7_n148 ) , .ZN( u0_u12_u7_n169 ) );
  INV_X1 u0_u12_u7_U34 (.A( u0_u12_u7_n127 ) , .ZN( u0_u12_u7_n179 ) );
  NOR2_X1 u0_u12_u7_U35 (.ZN( u0_u12_u7_n101 ) , .A2( u0_u12_u7_n150 ) , .A1( u0_u12_u7_n156 ) );
  AOI211_X1 u0_u12_u7_U36 (.B( u0_u12_u7_n154 ) , .A( u0_u12_u7_n155 ) , .C1( u0_u12_u7_n156 ) , .ZN( u0_u12_u7_n157 ) , .C2( u0_u12_u7_n172 ) );
  INV_X1 u0_u12_u7_U37 (.A( u0_u12_u7_n153 ) , .ZN( u0_u12_u7_n172 ) );
  AOI211_X1 u0_u12_u7_U38 (.B( u0_u12_u7_n139 ) , .A( u0_u12_u7_n140 ) , .C2( u0_u12_u7_n141 ) , .ZN( u0_u12_u7_n142 ) , .C1( u0_u12_u7_n156 ) );
  NAND4_X1 u0_u12_u7_U39 (.A3( u0_u12_u7_n127 ) , .A2( u0_u12_u7_n128 ) , .A1( u0_u12_u7_n129 ) , .ZN( u0_u12_u7_n141 ) , .A4( u0_u12_u7_n147 ) );
  INV_X1 u0_u12_u7_U4 (.A( u0_u12_u7_n111 ) , .ZN( u0_u12_u7_n170 ) );
  AOI21_X1 u0_u12_u7_U40 (.A( u0_u12_u7_n137 ) , .B1( u0_u12_u7_n138 ) , .ZN( u0_u12_u7_n139 ) , .B2( u0_u12_u7_n146 ) );
  OAI22_X1 u0_u12_u7_U41 (.B1( u0_u12_u7_n136 ) , .ZN( u0_u12_u7_n140 ) , .A1( u0_u12_u7_n153 ) , .B2( u0_u12_u7_n162 ) , .A2( u0_u12_u7_n164 ) );
  AOI21_X1 u0_u12_u7_U42 (.ZN( u0_u12_u7_n123 ) , .B1( u0_u12_u7_n165 ) , .B2( u0_u12_u7_n177 ) , .A( u0_u12_u7_n97 ) );
  AOI21_X1 u0_u12_u7_U43 (.B2( u0_u12_u7_n113 ) , .B1( u0_u12_u7_n124 ) , .A( u0_u12_u7_n125 ) , .ZN( u0_u12_u7_n97 ) );
  INV_X1 u0_u12_u7_U44 (.A( u0_u12_u7_n125 ) , .ZN( u0_u12_u7_n161 ) );
  INV_X1 u0_u12_u7_U45 (.A( u0_u12_u7_n152 ) , .ZN( u0_u12_u7_n162 ) );
  AOI22_X1 u0_u12_u7_U46 (.A2( u0_u12_u7_n114 ) , .ZN( u0_u12_u7_n119 ) , .B1( u0_u12_u7_n130 ) , .A1( u0_u12_u7_n156 ) , .B2( u0_u12_u7_n165 ) );
  NAND2_X1 u0_u12_u7_U47 (.A2( u0_u12_u7_n112 ) , .ZN( u0_u12_u7_n114 ) , .A1( u0_u12_u7_n175 ) );
  AND2_X1 u0_u12_u7_U48 (.ZN( u0_u12_u7_n145 ) , .A2( u0_u12_u7_n98 ) , .A1( u0_u12_u7_n99 ) );
  NOR2_X1 u0_u12_u7_U49 (.ZN( u0_u12_u7_n137 ) , .A1( u0_u12_u7_n150 ) , .A2( u0_u12_u7_n161 ) );
  INV_X1 u0_u12_u7_U5 (.A( u0_u12_u7_n149 ) , .ZN( u0_u12_u7_n175 ) );
  AOI21_X1 u0_u12_u7_U50 (.ZN( u0_u12_u7_n105 ) , .B2( u0_u12_u7_n110 ) , .A( u0_u12_u7_n125 ) , .B1( u0_u12_u7_n147 ) );
  NAND2_X1 u0_u12_u7_U51 (.ZN( u0_u12_u7_n146 ) , .A1( u0_u12_u7_n95 ) , .A2( u0_u12_u7_n98 ) );
  NAND2_X1 u0_u12_u7_U52 (.A2( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n147 ) , .A1( u0_u12_u7_n93 ) );
  NAND2_X1 u0_u12_u7_U53 (.A1( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n127 ) , .A2( u0_u12_u7_n99 ) );
  OR2_X1 u0_u12_u7_U54 (.ZN( u0_u12_u7_n126 ) , .A2( u0_u12_u7_n152 ) , .A1( u0_u12_u7_n156 ) );
  NAND2_X1 u0_u12_u7_U55 (.A2( u0_u12_u7_n102 ) , .A1( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n133 ) );
  NAND2_X1 u0_u12_u7_U56 (.ZN( u0_u12_u7_n112 ) , .A2( u0_u12_u7_n96 ) , .A1( u0_u12_u7_n99 ) );
  NAND2_X1 u0_u12_u7_U57 (.A2( u0_u12_u7_n102 ) , .ZN( u0_u12_u7_n128 ) , .A1( u0_u12_u7_n98 ) );
  NAND2_X1 u0_u12_u7_U58 (.A1( u0_u12_u7_n100 ) , .ZN( u0_u12_u7_n113 ) , .A2( u0_u12_u7_n93 ) );
  NAND2_X1 u0_u12_u7_U59 (.A2( u0_u12_u7_n102 ) , .ZN( u0_u12_u7_n124 ) , .A1( u0_u12_u7_n96 ) );
  INV_X1 u0_u12_u7_U6 (.A( u0_u12_u7_n154 ) , .ZN( u0_u12_u7_n178 ) );
  NAND2_X1 u0_u12_u7_U60 (.ZN( u0_u12_u7_n110 ) , .A1( u0_u12_u7_n95 ) , .A2( u0_u12_u7_n96 ) );
  INV_X1 u0_u12_u7_U61 (.A( u0_u12_u7_n150 ) , .ZN( u0_u12_u7_n164 ) );
  AND2_X1 u0_u12_u7_U62 (.ZN( u0_u12_u7_n134 ) , .A1( u0_u12_u7_n93 ) , .A2( u0_u12_u7_n98 ) );
  NAND2_X1 u0_u12_u7_U63 (.A1( u0_u12_u7_n100 ) , .A2( u0_u12_u7_n102 ) , .ZN( u0_u12_u7_n129 ) );
  NAND2_X1 u0_u12_u7_U64 (.A2( u0_u12_u7_n103 ) , .ZN( u0_u12_u7_n131 ) , .A1( u0_u12_u7_n95 ) );
  NAND2_X1 u0_u12_u7_U65 (.A1( u0_u12_u7_n100 ) , .ZN( u0_u12_u7_n138 ) , .A2( u0_u12_u7_n99 ) );
  NAND2_X1 u0_u12_u7_U66 (.ZN( u0_u12_u7_n132 ) , .A1( u0_u12_u7_n93 ) , .A2( u0_u12_u7_n96 ) );
  NAND2_X1 u0_u12_u7_U67 (.A1( u0_u12_u7_n100 ) , .ZN( u0_u12_u7_n148 ) , .A2( u0_u12_u7_n95 ) );
  NOR2_X1 u0_u12_u7_U68 (.A2( u0_u12_X_47 ) , .ZN( u0_u12_u7_n150 ) , .A1( u0_u12_u7_n163 ) );
  NOR2_X1 u0_u12_u7_U69 (.A2( u0_u12_X_43 ) , .A1( u0_u12_X_44 ) , .ZN( u0_u12_u7_n103 ) );
  AOI211_X1 u0_u12_u7_U7 (.ZN( u0_u12_u7_n116 ) , .A( u0_u12_u7_n155 ) , .C1( u0_u12_u7_n161 ) , .C2( u0_u12_u7_n171 ) , .B( u0_u12_u7_n94 ) );
  NOR2_X1 u0_u12_u7_U70 (.A2( u0_u12_X_48 ) , .A1( u0_u12_u7_n166 ) , .ZN( u0_u12_u7_n95 ) );
  NOR2_X1 u0_u12_u7_U71 (.A2( u0_u12_X_45 ) , .A1( u0_u12_X_48 ) , .ZN( u0_u12_u7_n99 ) );
  NOR2_X1 u0_u12_u7_U72 (.A2( u0_u12_X_44 ) , .A1( u0_u12_u7_n167 ) , .ZN( u0_u12_u7_n98 ) );
  NOR2_X1 u0_u12_u7_U73 (.A2( u0_u12_X_46 ) , .A1( u0_u12_X_47 ) , .ZN( u0_u12_u7_n152 ) );
  AND2_X1 u0_u12_u7_U74 (.A1( u0_u12_X_47 ) , .ZN( u0_u12_u7_n156 ) , .A2( u0_u12_u7_n163 ) );
  NAND2_X1 u0_u12_u7_U75 (.A2( u0_u12_X_46 ) , .A1( u0_u12_X_47 ) , .ZN( u0_u12_u7_n125 ) );
  AND2_X1 u0_u12_u7_U76 (.A2( u0_u12_X_45 ) , .A1( u0_u12_X_48 ) , .ZN( u0_u12_u7_n102 ) );
  AND2_X1 u0_u12_u7_U77 (.A2( u0_u12_X_43 ) , .A1( u0_u12_X_44 ) , .ZN( u0_u12_u7_n96 ) );
  AND2_X1 u0_u12_u7_U78 (.A1( u0_u12_X_44 ) , .ZN( u0_u12_u7_n100 ) , .A2( u0_u12_u7_n167 ) );
  AND2_X1 u0_u12_u7_U79 (.A1( u0_u12_X_48 ) , .A2( u0_u12_u7_n166 ) , .ZN( u0_u12_u7_n93 ) );
  OAI222_X1 u0_u12_u7_U8 (.C2( u0_u12_u7_n101 ) , .B2( u0_u12_u7_n111 ) , .A1( u0_u12_u7_n113 ) , .C1( u0_u12_u7_n146 ) , .A2( u0_u12_u7_n162 ) , .B1( u0_u12_u7_n164 ) , .ZN( u0_u12_u7_n94 ) );
  INV_X1 u0_u12_u7_U80 (.A( u0_u12_X_46 ) , .ZN( u0_u12_u7_n163 ) );
  INV_X1 u0_u12_u7_U81 (.A( u0_u12_X_43 ) , .ZN( u0_u12_u7_n167 ) );
  INV_X1 u0_u12_u7_U82 (.A( u0_u12_X_45 ) , .ZN( u0_u12_u7_n166 ) );
  NAND4_X1 u0_u12_u7_U83 (.ZN( u0_out12_27 ) , .A4( u0_u12_u7_n118 ) , .A3( u0_u12_u7_n119 ) , .A2( u0_u12_u7_n120 ) , .A1( u0_u12_u7_n121 ) );
  OAI21_X1 u0_u12_u7_U84 (.ZN( u0_u12_u7_n121 ) , .B2( u0_u12_u7_n145 ) , .A( u0_u12_u7_n150 ) , .B1( u0_u12_u7_n174 ) );
  OAI21_X1 u0_u12_u7_U85 (.ZN( u0_u12_u7_n120 ) , .A( u0_u12_u7_n161 ) , .B2( u0_u12_u7_n170 ) , .B1( u0_u12_u7_n179 ) );
  NAND4_X1 u0_u12_u7_U86 (.ZN( u0_out12_21 ) , .A4( u0_u12_u7_n157 ) , .A3( u0_u12_u7_n158 ) , .A2( u0_u12_u7_n159 ) , .A1( u0_u12_u7_n160 ) );
  OAI21_X1 u0_u12_u7_U87 (.B1( u0_u12_u7_n145 ) , .ZN( u0_u12_u7_n160 ) , .A( u0_u12_u7_n161 ) , .B2( u0_u12_u7_n177 ) );
  AOI22_X1 u0_u12_u7_U88 (.B2( u0_u12_u7_n149 ) , .B1( u0_u12_u7_n150 ) , .A2( u0_u12_u7_n151 ) , .A1( u0_u12_u7_n152 ) , .ZN( u0_u12_u7_n158 ) );
  NAND4_X1 u0_u12_u7_U89 (.ZN( u0_out12_15 ) , .A4( u0_u12_u7_n142 ) , .A3( u0_u12_u7_n143 ) , .A2( u0_u12_u7_n144 ) , .A1( u0_u12_u7_n178 ) );
  OAI221_X1 u0_u12_u7_U9 (.C1( u0_u12_u7_n101 ) , .C2( u0_u12_u7_n147 ) , .ZN( u0_u12_u7_n155 ) , .B2( u0_u12_u7_n162 ) , .A( u0_u12_u7_n91 ) , .B1( u0_u12_u7_n92 ) );
  OR2_X1 u0_u12_u7_U90 (.A2( u0_u12_u7_n125 ) , .A1( u0_u12_u7_n129 ) , .ZN( u0_u12_u7_n144 ) );
  AOI22_X1 u0_u12_u7_U91 (.A2( u0_u12_u7_n126 ) , .ZN( u0_u12_u7_n143 ) , .B2( u0_u12_u7_n165 ) , .B1( u0_u12_u7_n173 ) , .A1( u0_u12_u7_n174 ) );
  NAND4_X1 u0_u12_u7_U92 (.ZN( u0_out12_5 ) , .A4( u0_u12_u7_n108 ) , .A3( u0_u12_u7_n109 ) , .A1( u0_u12_u7_n116 ) , .A2( u0_u12_u7_n123 ) );
  AOI22_X1 u0_u12_u7_U93 (.ZN( u0_u12_u7_n109 ) , .A2( u0_u12_u7_n126 ) , .B2( u0_u12_u7_n145 ) , .B1( u0_u12_u7_n156 ) , .A1( u0_u12_u7_n171 ) );
  NOR4_X1 u0_u12_u7_U94 (.A4( u0_u12_u7_n104 ) , .A3( u0_u12_u7_n105 ) , .A2( u0_u12_u7_n106 ) , .A1( u0_u12_u7_n107 ) , .ZN( u0_u12_u7_n108 ) );
  NAND3_X1 u0_u12_u7_U95 (.A3( u0_u12_u7_n146 ) , .A2( u0_u12_u7_n147 ) , .A1( u0_u12_u7_n148 ) , .ZN( u0_u12_u7_n151 ) );
  NAND3_X1 u0_u12_u7_U96 (.A3( u0_u12_u7_n131 ) , .A2( u0_u12_u7_n132 ) , .A1( u0_u12_u7_n133 ) , .ZN( u0_u12_u7_n135 ) );
  OAI22_X1 u0_uk_U110 (.ZN( u0_K12_41 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n144 ) , .B1( u0_uk_n148 ) , .B2( u0_uk_n153 ) );
  OAI22_X1 u0_uk_U113 (.ZN( u0_K13_47 ) , .B2( u0_uk_n106 ) , .B1( u0_uk_n252 ) , .A2( u0_uk_n96 ) , .A1( u0_uk_n99 ) );
  INV_X1 u0_uk_U1131 (.ZN( u0_K12_42 ) , .A( u0_uk_n966 ) );
  AOI22_X1 u0_uk_U1132 (.B2( u0_uk_K_r10_28 ) , .A2( u0_uk_K_r10_9 ) , .B1( u0_uk_n129 ) , .A1( u0_uk_n213 ) , .ZN( u0_uk_n966 ) );
  OAI22_X1 u0_uk_U114 (.ZN( u0_K12_47 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n152 ) , .B2( u0_uk_n179 ) );
  INV_X1 u0_uk_U1159 (.ZN( u0_K13_6 ) , .A( u0_uk_n940 ) );
  INV_X1 u0_uk_U167 (.ZN( u0_K12_30 ) , .A( u0_uk_n974 ) );
  AOI22_X1 u0_uk_U168 (.B2( u0_uk_K_r10_23 ) , .A2( u0_uk_K_r10_42 ) , .A1( u0_uk_n145 ) , .B1( u0_uk_n203 ) , .ZN( u0_uk_n974 ) );
  INV_X1 u0_uk_U190 (.ZN( u0_K11_30 ) , .A( u0_uk_n993 ) );
  AOI22_X1 u0_uk_U191 (.B2( u0_uk_K_r9_1 ) , .A2( u0_uk_K_r9_9 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n163 ) , .ZN( u0_uk_n993 ) );
  OAI21_X1 u0_uk_U216 (.ZN( u0_K12_31 ) , .B2( u0_uk_n173 ) , .B1( u0_uk_n250 ) , .A( u0_uk_n973 ) );
  NAND2_X1 u0_uk_U217 (.A1( u0_uk_K_r10_44 ) , .A2( u0_uk_n208 ) , .ZN( u0_uk_n973 ) );
  OAI22_X1 u0_uk_U255 (.ZN( u0_K13_44 ) , .B1( u0_uk_n110 ) , .A2( u0_uk_n119 ) , .B2( u0_uk_n134 ) , .A1( u0_uk_n191 ) );
  INV_X1 u0_uk_U258 (.ZN( u0_K12_44 ) , .A( u0_uk_n965 ) );
  AOI22_X1 u0_uk_U259 (.B2( u0_uk_K_r10_37 ) , .A2( u0_uk_K_r10_42 ) , .B1( u0_uk_n145 ) , .A1( u0_uk_n161 ) , .ZN( u0_uk_n965 ) );
  OAI21_X1 u0_uk_U308 (.ZN( u0_K11_26 ) , .B2( u0_uk_n193 ) , .B1( u0_uk_n93 ) , .A( u0_uk_n995 ) );
  NAND2_X1 u0_uk_U309 (.A1( u0_uk_K_r9_35 ) , .A2( u0_uk_n92 ) , .ZN( u0_uk_n995 ) );
  OAI22_X1 u0_uk_U316 (.ZN( u0_K12_26 ) , .B2( u0_uk_n168 ) , .A2( u0_uk_n178 ) , .B1( u0_uk_n182 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U322 (.ZN( u0_K12_46 ) , .A2( u0_uk_n140 ) , .B2( u0_uk_n180 ) , .A1( u0_uk_n252 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U374 (.ZN( u0_K11_28 ) , .A1( u0_uk_n109 ) , .A2( u0_uk_n184 ) , .B2( u0_uk_n216 ) , .B1( u0_uk_n222 ) );
  OAI22_X1 u0_uk_U382 (.ZN( u0_K12_28 ) , .A1( u0_uk_n102 ) , .A2( u0_uk_n174 ) , .B2( u0_uk_n178 ) , .B1( u0_uk_n214 ) );
  OAI21_X1 u0_uk_U441 (.ZN( u0_K12_33 ) , .B1( u0_uk_n10 ) , .B2( u0_uk_n140 ) , .A( u0_uk_n971 ) );
  NAND2_X1 u0_uk_U442 (.A1( u0_uk_K_r10_14 ) , .A2( u0_uk_n118 ) , .ZN( u0_uk_n971 ) );
  OAI22_X1 u0_uk_U456 (.ZN( u0_K12_37 ) , .A2( u0_uk_n139 ) , .B2( u0_uk_n179 ) , .A1( u0_uk_n238 ) , .B1( u0_uk_n92 ) );
  OAI21_X1 u0_uk_U475 (.ZN( u0_K11_29 ) , .B1( u0_uk_n129 ) , .B2( u0_uk_n224 ) , .A( u0_uk_n994 ) );
  NAND2_X1 u0_uk_U476 (.A1( u0_uk_K_r9_0 ) , .A2( u0_uk_n60 ) , .ZN( u0_uk_n994 ) );
  OAI22_X1 u0_uk_U485 (.ZN( u0_K12_29 ) , .A2( u0_uk_n144 ) , .B2( u0_uk_n167 ) , .A1( u0_uk_n251 ) , .B1( u0_uk_n92 ) );
  OAI22_X1 u0_uk_U555 (.ZN( u0_K12_38 ) , .A1( u0_uk_n129 ) , .B1( u0_uk_n148 ) , .A2( u0_uk_n153 ) , .B2( u0_uk_n180 ) );
  OAI21_X1 u0_uk_U664 (.ZN( u0_K13_43 ) , .B1( u0_uk_n252 ) , .A( u0_uk_n943 ) , .B2( u0_uk_n96 ) );
  NAND2_X1 u0_uk_U665 (.A1( u0_uk_K_r11_29 ) , .A2( u0_uk_n207 ) , .ZN( u0_uk_n943 ) );
  OAI21_X1 u0_uk_U666 (.ZN( u0_K12_45 ) , .B2( u0_uk_n174 ) , .B1( u0_uk_n191 ) , .A( u0_uk_n964 ) );
  NAND2_X1 u0_uk_U667 (.A1( u0_uk_K_r10_43 ) , .A2( u0_uk_n203 ) , .ZN( u0_uk_n964 ) );
  OAI22_X1 u0_uk_U688 (.ZN( u0_K11_25 ) , .A2( u0_uk_n192 ) , .B2( u0_uk_n211 ) , .A1( u0_uk_n242 ) , .B1( u0_uk_n94 ) );
  OAI22_X1 u0_uk_U695 (.ZN( u0_K12_25 ) , .A1( u0_uk_n100 ) , .A2( u0_uk_n154 ) , .B2( u0_uk_n159 ) , .B1( u0_uk_n222 ) );
  INV_X1 u0_uk_U738 (.ZN( u0_K12_32 ) , .A( u0_uk_n972 ) );
  AOI22_X1 u0_uk_U739 (.B2( u0_uk_K_r10_23 ) , .A2( u0_uk_K_r10_28 ) , .A1( u0_uk_n251 ) , .B1( u0_uk_n60 ) , .ZN( u0_uk_n972 ) );
  OAI22_X1 u0_uk_U746 (.ZN( u0_K12_27 ) , .A2( u0_uk_n139 ) , .B2( u0_uk_n171 ) , .B1( u0_uk_n214 ) , .A1( u0_uk_n99 ) );
  OAI22_X1 u0_uk_U759 (.ZN( u0_K11_27 ) , .A1( u0_uk_n109 ) , .B1( u0_uk_n182 ) , .A2( u0_uk_n198 ) , .B2( u0_uk_n204 ) );
  OAI21_X1 u0_uk_U835 (.ZN( u0_K13_1 ) , .B2( u0_uk_n131 ) , .B1( u0_uk_n31 ) , .A( u0_uk_n952 ) );
  NAND2_X1 u0_uk_U836 (.A1( u0_uk_K_r11_25 ) , .A2( u0_uk_n11 ) , .ZN( u0_uk_n952 ) );
  OAI21_X1 u0_uk_U847 (.ZN( u0_K13_3 ) , .B2( u0_uk_n107 ) , .B1( u0_uk_n31 ) , .A( u0_uk_n944 ) );
  NAND2_X1 u0_uk_U848 (.A1( u0_uk_K_r11_4 ) , .A2( u0_uk_n129 ) , .ZN( u0_uk_n944 ) );
  INV_X1 u0_uk_U852 (.ZN( u0_K13_2 ) , .A( u0_uk_n946 ) );
  AOI22_X1 u0_uk_U853 (.B2( u0_uk_K_r11_26 ) , .A2( u0_uk_K_r11_46 ) , .A1( u0_uk_n10 ) , .B1( u0_uk_n163 ) , .ZN( u0_uk_n946 ) );
  AOI22_X1 u0_uk_U866 (.B2( u0_uk_K_r11_19 ) , .A2( u0_uk_K_r11_24 ) , .B1( u0_uk_n142 ) , .A1( u0_uk_n217 ) , .ZN( u0_uk_n940 ) );
  OAI22_X1 u0_uk_U888 (.ZN( u0_K12_43 ) , .A2( u0_uk_n151 ) , .B2( u0_uk_n171 ) , .A1( u0_uk_n220 ) , .B1( u0_uk_n83 ) );
  OAI22_X1 u0_uk_U952 (.ZN( u0_K13_4 ) , .A1( u0_uk_n117 ) , .A2( u0_uk_n121 ) , .B2( u0_uk_n126 ) , .B1( u0_uk_n214 ) );
  INV_X1 u0_uk_U98 (.ZN( u0_K13_5 ) , .A( u0_uk_n941 ) );
  AOI22_X1 u0_uk_U99 (.B2( u0_uk_K_r11_48 ) , .A2( u0_uk_K_r11_53 ) , .B1( u0_uk_n141 ) , .A1( u0_uk_n220 ) , .ZN( u0_uk_n941 ) );
  XOR2_X1 u2_U100 (.B( u2_L12_27 ) , .Z( u2_N442 ) , .A( u2_out13_27 ) );
  XOR2_X1 u2_U107 (.B( u2_L12_21 ) , .Z( u2_N436 ) , .A( u2_out13_21 ) );
  XOR2_X1 u2_U113 (.B( u2_L12_15 ) , .Z( u2_N430 ) , .A( u2_out13_15 ) );
  XOR2_X1 u2_U114 (.B( u2_L0_12 ) , .Z( u2_N43 ) , .A( u2_out1_12 ) );
  XOR2_X1 u2_U124 (.B( u2_L12_5 ) , .Z( u2_N420 ) , .A( u2_out13_5 ) );
  XOR2_X1 u2_U125 (.B( u2_L0_11 ) , .Z( u2_N42 ) , .A( u2_out1_11 ) );
  XOR2_X1 u2_U13 (.Z( u2_N9 ) , .B( u2_desIn_r_12 ) , .A( u2_out0_10 ) );
  XOR2_X1 u2_U148 (.Z( u2_N4 ) , .B( u2_desIn_r_38 ) , .A( u2_out0_5 ) );
  XOR2_X1 u2_U167 (.B( u2_L10_31 ) , .Z( u2_N382 ) , .A( u2_out11_31 ) );
  XOR2_X1 u2_U170 (.B( u2_L0_7 ) , .Z( u2_N38 ) , .A( u2_out1_7 ) );
  XOR2_X1 u2_U171 (.B( u2_L10_28 ) , .Z( u2_N379 ) , .A( u2_out11_28 ) );
  XOR2_X1 u2_U176 (.B( u2_L10_23 ) , .Z( u2_N374 ) , .A( u2_out11_23 ) );
  XOR2_X1 u2_U182 (.B( u2_L10_18 ) , .Z( u2_N369 ) , .A( u2_out11_18 ) );
  XOR2_X1 u2_U183 (.B( u2_L10_17 ) , .Z( u2_N368 ) , .A( u2_out11_17 ) );
  XOR2_X1 u2_U187 (.B( u2_L10_13 ) , .Z( u2_N364 ) , .A( u2_out11_13 ) );
  XOR2_X1 u2_U191 (.B( u2_L10_9 ) , .Z( u2_N360 ) , .A( u2_out11_9 ) );
  XOR2_X1 u2_U199 (.B( u2_L10_2 ) , .Z( u2_N353 ) , .A( u2_out11_2 ) );
  XOR2_X1 u2_U203 (.B( u2_L0_4 ) , .Z( u2_N35 ) , .A( u2_out1_4 ) );
  XOR2_X1 u2_U237 (.B( u2_L8_32 ) , .Z( u2_N319 ) , .A( u2_out9_32 ) );
  XOR2_X1 u2_U240 (.B( u2_L8_29 ) , .Z( u2_N316 ) , .A( u2_out9_29 ) );
  XOR2_X1 u2_U247 (.Z( u2_N31 ) , .B( u2_desIn_r_56 ) , .A( u2_out0_32 ) );
  XOR2_X1 u2_U248 (.B( u2_L8_22 ) , .Z( u2_N309 ) , .A( u2_out9_22 ) );
  XOR2_X1 u2_U251 (.B( u2_L8_19 ) , .Z( u2_N306 ) , .A( u2_out9_19 ) );
  XOR2_X1 u2_U259 (.Z( u2_N3 ) , .B( u2_desIn_r_30 ) , .A( u2_out0_4 ) );
  XOR2_X1 u2_U260 (.B( u2_L8_12 ) , .Z( u2_N299 ) , .A( u2_out9_12 ) );
  XOR2_X1 u2_U261 (.B( u2_L8_11 ) , .Z( u2_N298 ) , .A( u2_out9_11 ) );
  XOR2_X1 u2_U265 (.B( u2_L8_7 ) , .Z( u2_N294 ) , .A( u2_out9_7 ) );
  XOR2_X1 u2_U268 (.B( u2_L8_4 ) , .Z( u2_N291 ) , .A( u2_out9_4 ) );
  XOR2_X1 u2_U279 (.B( u2_L7_26 ) , .Z( u2_N281 ) , .A( u2_out8_26 ) );
  XOR2_X1 u2_U280 (.B( u2_L7_25 ) , .Z( u2_N280 ) , .A( u2_out8_25 ) );
  XOR2_X1 u2_U281 (.Z( u2_N28 ) , .B( u2_desIn_r_32 ) , .A( u2_out0_29 ) );
  XOR2_X1 u2_U286 (.B( u2_L7_20 ) , .Z( u2_N275 ) , .A( u2_out8_20 ) );
  XOR2_X1 u2_U293 (.B( u2_L7_14 ) , .Z( u2_N269 ) , .A( u2_out8_14 ) );
  XOR2_X1 u2_U297 (.B( u2_L7_10 ) , .Z( u2_N265 ) , .A( u2_out8_10 ) );
  XOR2_X1 u2_U299 (.B( u2_L7_8 ) , .Z( u2_N263 ) , .A( u2_out8_8 ) );
  XOR2_X1 u2_U303 (.Z( u2_N26 ) , .B( u2_desIn_r_16 ) , .A( u2_out0_27 ) );
  XOR2_X1 u2_U305 (.B( u2_L7_3 ) , .Z( u2_N258 ) , .A( u2_out8_3 ) );
  XOR2_X1 u2_U307 (.B( u2_L7_1 ) , .Z( u2_N256 ) , .A( u2_out8_1 ) );
  XOR2_X1 u2_U309 (.B( u2_L6_31 ) , .Z( u2_N254 ) , .A( u2_out7_31 ) );
  XOR2_X1 u2_U310 (.B( u2_L6_30 ) , .Z( u2_N253 ) , .A( u2_out7_30 ) );
  XOR2_X1 u2_U314 (.Z( u2_N25 ) , .B( u2_desIn_r_8 ) , .A( u2_out0_26 ) );
  XOR2_X1 u2_U317 (.B( u2_L6_24 ) , .Z( u2_N247 ) , .A( u2_out7_24 ) );
  XOR2_X1 u2_U318 (.B( u2_L6_23 ) , .Z( u2_N246 ) , .A( u2_out7_23 ) );
  XOR2_X1 u2_U324 (.B( u2_L6_17 ) , .Z( u2_N240 ) , .A( u2_out7_17 ) );
  XOR2_X1 u2_U325 (.Z( u2_N24 ) , .B( u2_desIn_r_0 ) , .A( u2_out0_25 ) );
  XOR2_X1 u2_U326 (.B( u2_L6_16 ) , .Z( u2_N239 ) , .A( u2_out7_16 ) );
  XOR2_X1 u2_U333 (.B( u2_L6_9 ) , .Z( u2_N232 ) , .A( u2_out7_9 ) );
  XOR2_X1 u2_U337 (.B( u2_L6_6 ) , .Z( u2_N229 ) , .A( u2_out7_6 ) );
  XOR2_X1 u2_U35 (.Z( u2_N7 ) , .B( u2_desIn_r_62 ) , .A( u2_out0_8 ) );
  XOR2_X1 u2_U358 (.Z( u2_N21 ) , .B( u2_desIn_r_42 ) , .A( u2_out0_22 ) );
  XOR2_X1 u2_U369 (.Z( u2_N20 ) , .B( u2_desIn_r_34 ) , .A( u2_out0_21 ) );
  XOR2_X1 u2_U370 (.Z( u2_N2 ) , .B( u2_desIn_r_22 ) , .A( u2_out0_3 ) );
  XOR2_X1 u2_U381 (.Z( u2_N19 ) , .B( u2_desIn_r_26 ) , .A( u2_out0_20 ) );
  XOR2_X1 u2_U392 (.Z( u2_N18 ) , .B( u2_desIn_r_18 ) , .A( u2_out0_19 ) );
  XOR2_X1 u2_U416 (.B( u2_L3_31 ) , .Z( u2_N158 ) , .A( u2_out4_31 ) );
  XOR2_X1 u2_U417 (.B( u2_L3_30 ) , .Z( u2_N157 ) , .A( u2_out4_30 ) );
  XOR2_X1 u2_U419 (.B( u2_L3_28 ) , .Z( u2_N155 ) , .A( u2_out4_28 ) );
  XOR2_X1 u2_U42 (.B( u2_L0_32 ) , .Z( u2_N63 ) , .A( u2_out1_32 ) );
  XOR2_X1 u2_U421 (.B( u2_L3_26 ) , .Z( u2_N153 ) , .A( u2_out4_26 ) );
  XOR2_X1 u2_U422 (.B( u2_L3_25 ) , .Z( u2_N152 ) , .A( u2_out4_25 ) );
  XOR2_X1 u2_U423 (.B( u2_L3_24 ) , .Z( u2_N151 ) , .A( u2_out4_24 ) );
  XOR2_X1 u2_U424 (.B( u2_L3_23 ) , .Z( u2_N150 ) , .A( u2_out4_23 ) );
  XOR2_X1 u2_U428 (.B( u2_L3_20 ) , .Z( u2_N147 ) , .A( u2_out4_20 ) );
  XOR2_X1 u2_U430 (.B( u2_L3_18 ) , .Z( u2_N145 ) , .A( u2_out4_18 ) );
  XOR2_X1 u2_U431 (.B( u2_L3_17 ) , .Z( u2_N144 ) , .A( u2_out4_17 ) );
  XOR2_X1 u2_U432 (.B( u2_L3_16 ) , .Z( u2_N143 ) , .A( u2_out4_16 ) );
  XOR2_X1 u2_U434 (.B( u2_L3_14 ) , .Z( u2_N141 ) , .A( u2_out4_14 ) );
  XOR2_X1 u2_U435 (.B( u2_L3_13 ) , .Z( u2_N140 ) , .A( u2_out4_13 ) );
  XOR2_X1 u2_U436 (.Z( u2_N14 ) , .B( u2_desIn_r_52 ) , .A( u2_out0_15 ) );
  XOR2_X1 u2_U439 (.B( u2_L3_10 ) , .Z( u2_N137 ) , .A( u2_out4_10 ) );
  XOR2_X1 u2_U440 (.B( u2_L3_9 ) , .Z( u2_N136 ) , .A( u2_out4_9 ) );
  XOR2_X1 u2_U441 (.B( u2_L3_8 ) , .Z( u2_N135 ) , .A( u2_out4_8 ) );
  XOR2_X1 u2_U443 (.B( u2_L3_6 ) , .Z( u2_N133 ) , .A( u2_out4_6 ) );
  XOR2_X1 u2_U446 (.B( u2_L3_3 ) , .Z( u2_N130 ) , .A( u2_out4_3 ) );
  XOR2_X1 u2_U447 (.Z( u2_N13 ) , .B( u2_desIn_r_44 ) , .A( u2_out0_14 ) );
  XOR2_X1 u2_U448 (.B( u2_L3_2 ) , .Z( u2_N129 ) , .A( u2_out4_2 ) );
  XOR2_X1 u2_U449 (.B( u2_L3_1 ) , .Z( u2_N128 ) , .A( u2_out4_1 ) );
  XOR2_X1 u2_U45 (.B( u2_L0_29 ) , .Z( u2_N60 ) , .A( u2_out1_29 ) );
  XOR2_X1 u2_U46 (.Z( u2_N6 ) , .B( u2_desIn_r_54 ) , .A( u2_out0_7 ) );
  XOR2_X1 u2_U469 (.Z( u2_N11 ) , .B( u2_desIn_r_28 ) , .A( u2_out0_12 ) );
  XOR2_X1 u2_U480 (.Z( u2_N10 ) , .B( u2_desIn_r_20 ) , .A( u2_out0_11 ) );
  XOR2_X1 u2_U482 (.Z( u2_N0 ) , .B( u2_desIn_r_6 ) , .A( u2_out0_1 ) );
  XOR2_X1 u2_U53 (.B( u2_L0_22 ) , .Z( u2_N53 ) , .A( u2_out1_22 ) );
  XOR2_X1 u2_U56 (.B( u2_L0_19 ) , .Z( u2_N50 ) , .A( u2_out1_19 ) );
  XOR2_X1 u2_u0_U10 (.B( u2_K1_45 ) , .A( u2_desIn_r_41 ) , .Z( u2_u0_X_45 ) );
  XOR2_X1 u2_u0_U11 (.B( u2_K1_44 ) , .A( u2_desIn_r_33 ) , .Z( u2_u0_X_44 ) );
  XOR2_X1 u2_u0_U12 (.B( u2_K1_43 ) , .A( u2_desIn_r_25 ) , .Z( u2_u0_X_43 ) );
  XOR2_X1 u2_u0_U13 (.B( u2_K1_42 ) , .A( u2_desIn_r_33 ) , .Z( u2_u0_X_42 ) );
  XOR2_X1 u2_u0_U14 (.B( u2_K1_41 ) , .A( u2_desIn_r_25 ) , .Z( u2_u0_X_41 ) );
  XOR2_X1 u2_u0_U15 (.B( u2_K1_40 ) , .A( u2_desIn_r_17 ) , .Z( u2_u0_X_40 ) );
  XOR2_X1 u2_u0_U17 (.B( u2_K1_39 ) , .A( u2_desIn_r_9 ) , .Z( u2_u0_X_39 ) );
  XOR2_X1 u2_u0_U18 (.B( u2_K1_38 ) , .A( u2_desIn_r_1 ) , .Z( u2_u0_X_38 ) );
  XOR2_X1 u2_u0_U19 (.B( u2_K1_37 ) , .A( u2_desIn_r_59 ) , .Z( u2_u0_X_37 ) );
  XOR2_X1 u2_u0_U20 (.B( u2_K1_36 ) , .A( u2_desIn_r_1 ) , .Z( u2_u0_X_36 ) );
  XOR2_X1 u2_u0_U21 (.B( u2_K1_35 ) , .A( u2_desIn_r_59 ) , .Z( u2_u0_X_35 ) );
  XOR2_X1 u2_u0_U22 (.B( u2_K1_34 ) , .A( u2_desIn_r_51 ) , .Z( u2_u0_X_34 ) );
  XOR2_X1 u2_u0_U23 (.B( u2_K1_33 ) , .A( u2_desIn_r_43 ) , .Z( u2_u0_X_33 ) );
  XOR2_X1 u2_u0_U24 (.B( u2_K1_32 ) , .A( u2_desIn_r_35 ) , .Z( u2_u0_X_32 ) );
  XOR2_X1 u2_u0_U25 (.B( u2_K1_31 ) , .A( u2_desIn_r_27 ) , .Z( u2_u0_X_31 ) );
  XOR2_X1 u2_u0_U26 (.B( u2_K1_30 ) , .A( u2_desIn_r_35 ) , .Z( u2_u0_X_30 ) );
  XOR2_X1 u2_u0_U28 (.B( u2_K1_29 ) , .A( u2_desIn_r_27 ) , .Z( u2_u0_X_29 ) );
  XOR2_X1 u2_u0_U29 (.B( u2_K1_28 ) , .A( u2_desIn_r_19 ) , .Z( u2_u0_X_28 ) );
  XOR2_X1 u2_u0_U30 (.B( u2_K1_27 ) , .A( u2_desIn_r_11 ) , .Z( u2_u0_X_27 ) );
  XOR2_X1 u2_u0_U31 (.B( u2_K1_26 ) , .A( u2_desIn_r_3 ) , .Z( u2_u0_X_26 ) );
  XOR2_X1 u2_u0_U32 (.B( u2_K1_25 ) , .A( u2_desIn_r_61 ) , .Z( u2_u0_X_25 ) );
  XOR2_X1 u2_u0_U33 (.B( u2_K1_24 ) , .A( u2_desIn_r_3 ) , .Z( u2_u0_X_24 ) );
  XOR2_X1 u2_u0_U34 (.B( u2_K1_23 ) , .A( u2_desIn_r_61 ) , .Z( u2_u0_X_23 ) );
  XOR2_X1 u2_u0_U35 (.B( u2_K1_22 ) , .A( u2_desIn_r_53 ) , .Z( u2_u0_X_22 ) );
  XOR2_X1 u2_u0_U36 (.B( u2_K1_21 ) , .A( u2_desIn_r_45 ) , .Z( u2_u0_X_21 ) );
  XOR2_X1 u2_u0_U37 (.B( u2_K1_20 ) , .A( u2_desIn_r_37 ) , .Z( u2_u0_X_20 ) );
  XOR2_X1 u2_u0_U38 (.B( u2_K1_1 ) , .A( u2_desIn_r_57 ) , .Z( u2_u0_X_1 ) );
  XOR2_X1 u2_u0_U39 (.B( u2_K1_19 ) , .A( u2_desIn_r_29 ) , .Z( u2_u0_X_19 ) );
  XOR2_X1 u2_u0_U7 (.B( u2_K1_48 ) , .A( u2_desIn_r_7 ) , .Z( u2_u0_X_48 ) );
  XOR2_X1 u2_u0_U8 (.B( u2_K1_47 ) , .A( u2_desIn_r_57 ) , .Z( u2_u0_X_47 ) );
  XOR2_X1 u2_u0_U9 (.B( u2_K1_46 ) , .A( u2_desIn_r_49 ) , .Z( u2_u0_X_46 ) );
  OAI211_X1 u2_u0_u3_U10 (.B( u2_u0_u3_n106 ) , .ZN( u2_u0_u3_n119 ) , .C2( u2_u0_u3_n128 ) , .C1( u2_u0_u3_n167 ) , .A( u2_u0_u3_n181 ) );
  AOI221_X1 u2_u0_u3_U11 (.C1( u2_u0_u3_n105 ) , .ZN( u2_u0_u3_n106 ) , .A( u2_u0_u3_n131 ) , .B2( u2_u0_u3_n132 ) , .C2( u2_u0_u3_n133 ) , .B1( u2_u0_u3_n169 ) );
  INV_X1 u2_u0_u3_U12 (.ZN( u2_u0_u3_n181 ) , .A( u2_u0_u3_n98 ) );
  NAND2_X1 u2_u0_u3_U13 (.ZN( u2_u0_u3_n105 ) , .A2( u2_u0_u3_n130 ) , .A1( u2_u0_u3_n155 ) );
  AOI22_X1 u2_u0_u3_U14 (.B1( u2_u0_u3_n115 ) , .A2( u2_u0_u3_n116 ) , .ZN( u2_u0_u3_n123 ) , .B2( u2_u0_u3_n133 ) , .A1( u2_u0_u3_n169 ) );
  NAND2_X1 u2_u0_u3_U15 (.ZN( u2_u0_u3_n116 ) , .A2( u2_u0_u3_n151 ) , .A1( u2_u0_u3_n182 ) );
  NOR2_X1 u2_u0_u3_U16 (.ZN( u2_u0_u3_n126 ) , .A2( u2_u0_u3_n150 ) , .A1( u2_u0_u3_n164 ) );
  AOI21_X1 u2_u0_u3_U17 (.ZN( u2_u0_u3_n112 ) , .B2( u2_u0_u3_n146 ) , .B1( u2_u0_u3_n155 ) , .A( u2_u0_u3_n167 ) );
  NAND2_X1 u2_u0_u3_U18 (.A1( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n142 ) , .A2( u2_u0_u3_n164 ) );
  NAND2_X1 u2_u0_u3_U19 (.ZN( u2_u0_u3_n132 ) , .A2( u2_u0_u3_n152 ) , .A1( u2_u0_u3_n156 ) );
  INV_X1 u2_u0_u3_U20 (.A( u2_u0_u3_n133 ) , .ZN( u2_u0_u3_n165 ) );
  AND2_X1 u2_u0_u3_U21 (.A2( u2_u0_u3_n113 ) , .A1( u2_u0_u3_n114 ) , .ZN( u2_u0_u3_n151 ) );
  INV_X1 u2_u0_u3_U22 (.A( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n170 ) );
  NAND2_X1 u2_u0_u3_U23 (.A1( u2_u0_u3_n107 ) , .A2( u2_u0_u3_n108 ) , .ZN( u2_u0_u3_n140 ) );
  NAND2_X1 u2_u0_u3_U24 (.ZN( u2_u0_u3_n117 ) , .A1( u2_u0_u3_n124 ) , .A2( u2_u0_u3_n148 ) );
  INV_X1 u2_u0_u3_U25 (.A( u2_u0_u3_n128 ) , .ZN( u2_u0_u3_n176 ) );
  INV_X1 u2_u0_u3_U26 (.A( u2_u0_u3_n155 ) , .ZN( u2_u0_u3_n174 ) );
  INV_X1 u2_u0_u3_U27 (.A( u2_u0_u3_n130 ) , .ZN( u2_u0_u3_n177 ) );
  INV_X1 u2_u0_u3_U28 (.A( u2_u0_u3_n139 ) , .ZN( u2_u0_u3_n185 ) );
  NOR2_X1 u2_u0_u3_U29 (.ZN( u2_u0_u3_n135 ) , .A2( u2_u0_u3_n141 ) , .A1( u2_u0_u3_n169 ) );
  INV_X1 u2_u0_u3_U3 (.A( u2_u0_u3_n140 ) , .ZN( u2_u0_u3_n182 ) );
  OAI222_X1 u2_u0_u3_U30 (.C2( u2_u0_u3_n107 ) , .A2( u2_u0_u3_n108 ) , .B1( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n138 ) , .B2( u2_u0_u3_n146 ) , .C1( u2_u0_u3_n154 ) , .A1( u2_u0_u3_n164 ) );
  NOR4_X1 u2_u0_u3_U31 (.A4( u2_u0_u3_n157 ) , .A3( u2_u0_u3_n158 ) , .A2( u2_u0_u3_n159 ) , .A1( u2_u0_u3_n160 ) , .ZN( u2_u0_u3_n161 ) );
  AOI21_X1 u2_u0_u3_U32 (.B2( u2_u0_u3_n152 ) , .B1( u2_u0_u3_n153 ) , .ZN( u2_u0_u3_n158 ) , .A( u2_u0_u3_n164 ) );
  AOI21_X1 u2_u0_u3_U33 (.A( u2_u0_u3_n154 ) , .B2( u2_u0_u3_n155 ) , .B1( u2_u0_u3_n156 ) , .ZN( u2_u0_u3_n157 ) );
  AOI21_X1 u2_u0_u3_U34 (.A( u2_u0_u3_n149 ) , .B2( u2_u0_u3_n150 ) , .B1( u2_u0_u3_n151 ) , .ZN( u2_u0_u3_n159 ) );
  AOI211_X1 u2_u0_u3_U35 (.ZN( u2_u0_u3_n109 ) , .A( u2_u0_u3_n119 ) , .C2( u2_u0_u3_n129 ) , .B( u2_u0_u3_n138 ) , .C1( u2_u0_u3_n141 ) );
  AOI211_X1 u2_u0_u3_U36 (.B( u2_u0_u3_n119 ) , .A( u2_u0_u3_n120 ) , .C2( u2_u0_u3_n121 ) , .ZN( u2_u0_u3_n122 ) , .C1( u2_u0_u3_n179 ) );
  INV_X1 u2_u0_u3_U37 (.A( u2_u0_u3_n156 ) , .ZN( u2_u0_u3_n179 ) );
  OAI22_X1 u2_u0_u3_U38 (.B1( u2_u0_u3_n118 ) , .ZN( u2_u0_u3_n120 ) , .A1( u2_u0_u3_n135 ) , .B2( u2_u0_u3_n154 ) , .A2( u2_u0_u3_n178 ) );
  AND3_X1 u2_u0_u3_U39 (.ZN( u2_u0_u3_n118 ) , .A2( u2_u0_u3_n124 ) , .A1( u2_u0_u3_n144 ) , .A3( u2_u0_u3_n152 ) );
  INV_X1 u2_u0_u3_U4 (.A( u2_u0_u3_n129 ) , .ZN( u2_u0_u3_n183 ) );
  INV_X1 u2_u0_u3_U40 (.A( u2_u0_u3_n121 ) , .ZN( u2_u0_u3_n164 ) );
  OAI211_X1 u2_u0_u3_U41 (.B( u2_u0_u3_n127 ) , .ZN( u2_u0_u3_n139 ) , .C1( u2_u0_u3_n150 ) , .C2( u2_u0_u3_n154 ) , .A( u2_u0_u3_n184 ) );
  INV_X1 u2_u0_u3_U42 (.A( u2_u0_u3_n125 ) , .ZN( u2_u0_u3_n184 ) );
  AOI221_X1 u2_u0_u3_U43 (.A( u2_u0_u3_n126 ) , .ZN( u2_u0_u3_n127 ) , .C2( u2_u0_u3_n132 ) , .C1( u2_u0_u3_n169 ) , .B2( u2_u0_u3_n170 ) , .B1( u2_u0_u3_n174 ) );
  OAI22_X1 u2_u0_u3_U44 (.A1( u2_u0_u3_n124 ) , .ZN( u2_u0_u3_n125 ) , .B2( u2_u0_u3_n145 ) , .A2( u2_u0_u3_n165 ) , .B1( u2_u0_u3_n167 ) );
  NAND2_X1 u2_u0_u3_U45 (.A1( u2_u0_u3_n103 ) , .ZN( u2_u0_u3_n150 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U46 (.A2( u2_u0_u3_n102 ) , .ZN( u2_u0_u3_n155 ) , .A1( u2_u0_u3_n97 ) );
  NAND2_X1 u2_u0_u3_U47 (.ZN( u2_u0_u3_n133 ) , .A1( u2_u0_u3_n154 ) , .A2( u2_u0_u3_n164 ) );
  NOR2_X1 u2_u0_u3_U48 (.A1( u2_u0_u3_n113 ) , .ZN( u2_u0_u3_n131 ) , .A2( u2_u0_u3_n154 ) );
  AOI21_X1 u2_u0_u3_U49 (.B2( u2_u0_u3_n114 ) , .B1( u2_u0_u3_n146 ) , .A( u2_u0_u3_n154 ) , .ZN( u2_u0_u3_n94 ) );
  INV_X1 u2_u0_u3_U5 (.A( u2_u0_u3_n117 ) , .ZN( u2_u0_u3_n178 ) );
  AOI21_X1 u2_u0_u3_U50 (.ZN( u2_u0_u3_n110 ) , .B2( u2_u0_u3_n142 ) , .B1( u2_u0_u3_n186 ) , .A( u2_u0_u3_n95 ) );
  INV_X1 u2_u0_u3_U51 (.A( u2_u0_u3_n145 ) , .ZN( u2_u0_u3_n186 ) );
  AOI21_X1 u2_u0_u3_U52 (.B1( u2_u0_u3_n124 ) , .A( u2_u0_u3_n149 ) , .B2( u2_u0_u3_n155 ) , .ZN( u2_u0_u3_n95 ) );
  INV_X1 u2_u0_u3_U53 (.A( u2_u0_u3_n141 ) , .ZN( u2_u0_u3_n167 ) );
  NAND2_X1 u2_u0_u3_U54 (.ZN( u2_u0_u3_n124 ) , .A1( u2_u0_u3_n96 ) , .A2( u2_u0_u3_n97 ) );
  NAND2_X1 u2_u0_u3_U55 (.A2( u2_u0_u3_n100 ) , .ZN( u2_u0_u3_n146 ) , .A1( u2_u0_u3_n96 ) );
  INV_X1 u2_u0_u3_U56 (.A( u2_u0_u3_n149 ) , .ZN( u2_u0_u3_n169 ) );
  NAND2_X1 u2_u0_u3_U57 (.A1( u2_u0_u3_n101 ) , .ZN( u2_u0_u3_n145 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U58 (.A1( u2_u0_u3_n100 ) , .ZN( u2_u0_u3_n156 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U59 (.A2( u2_u0_u3_n101 ) , .A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n148 ) );
  OAI22_X1 u2_u0_u3_U6 (.B2( u2_u0_u3_n147 ) , .A2( u2_u0_u3_n148 ) , .ZN( u2_u0_u3_n160 ) , .B1( u2_u0_u3_n165 ) , .A1( u2_u0_u3_n168 ) );
  NAND2_X1 u2_u0_u3_U60 (.A1( u2_u0_u3_n100 ) , .A2( u2_u0_u3_n102 ) , .ZN( u2_u0_u3_n128 ) );
  NAND2_X1 u2_u0_u3_U61 (.A2( u2_u0_u3_n101 ) , .A1( u2_u0_u3_n102 ) , .ZN( u2_u0_u3_n152 ) );
  NAND2_X1 u2_u0_u3_U62 (.A2( u2_u0_u3_n101 ) , .ZN( u2_u0_u3_n114 ) , .A1( u2_u0_u3_n96 ) );
  NAND2_X1 u2_u0_u3_U63 (.ZN( u2_u0_u3_n107 ) , .A1( u2_u0_u3_n97 ) , .A2( u2_u0_u3_n99 ) );
  NAND2_X1 u2_u0_u3_U64 (.A2( u2_u0_u3_n100 ) , .A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n113 ) );
  NAND2_X1 u2_u0_u3_U65 (.A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n153 ) , .A2( u2_u0_u3_n97 ) );
  NAND2_X1 u2_u0_u3_U66 (.A2( u2_u0_u3_n103 ) , .A1( u2_u0_u3_n104 ) , .ZN( u2_u0_u3_n130 ) );
  NAND2_X1 u2_u0_u3_U67 (.A2( u2_u0_u3_n103 ) , .ZN( u2_u0_u3_n144 ) , .A1( u2_u0_u3_n96 ) );
  NAND2_X1 u2_u0_u3_U68 (.A1( u2_u0_u3_n102 ) , .A2( u2_u0_u3_n103 ) , .ZN( u2_u0_u3_n108 ) );
  NOR2_X1 u2_u0_u3_U69 (.A2( u2_u0_X_19 ) , .A1( u2_u0_X_20 ) , .ZN( u2_u0_u3_n99 ) );
  AND3_X1 u2_u0_u3_U7 (.A3( u2_u0_u3_n144 ) , .A2( u2_u0_u3_n145 ) , .A1( u2_u0_u3_n146 ) , .ZN( u2_u0_u3_n147 ) );
  NOR2_X1 u2_u0_u3_U70 (.A2( u2_u0_X_21 ) , .A1( u2_u0_X_24 ) , .ZN( u2_u0_u3_n103 ) );
  NOR2_X1 u2_u0_u3_U71 (.A2( u2_u0_X_24 ) , .A1( u2_u0_u3_n171 ) , .ZN( u2_u0_u3_n97 ) );
  NOR2_X1 u2_u0_u3_U72 (.A2( u2_u0_X_23 ) , .ZN( u2_u0_u3_n141 ) , .A1( u2_u0_u3_n166 ) );
  NOR2_X1 u2_u0_u3_U73 (.A2( u2_u0_X_19 ) , .A1( u2_u0_u3_n172 ) , .ZN( u2_u0_u3_n96 ) );
  NAND2_X1 u2_u0_u3_U74 (.A1( u2_u0_X_22 ) , .A2( u2_u0_X_23 ) , .ZN( u2_u0_u3_n154 ) );
  NOR2_X1 u2_u0_u3_U75 (.A2( u2_u0_X_22 ) , .A1( u2_u0_X_23 ) , .ZN( u2_u0_u3_n121 ) );
  AND2_X1 u2_u0_u3_U76 (.A1( u2_u0_X_24 ) , .ZN( u2_u0_u3_n101 ) , .A2( u2_u0_u3_n171 ) );
  NAND2_X1 u2_u0_u3_U77 (.A1( u2_u0_X_23 ) , .ZN( u2_u0_u3_n149 ) , .A2( u2_u0_u3_n166 ) );
  AND2_X1 u2_u0_u3_U78 (.A1( u2_u0_X_19 ) , .ZN( u2_u0_u3_n102 ) , .A2( u2_u0_u3_n172 ) );
  AND2_X1 u2_u0_u3_U79 (.A1( u2_u0_X_21 ) , .A2( u2_u0_X_24 ) , .ZN( u2_u0_u3_n100 ) );
  INV_X1 u2_u0_u3_U8 (.A( u2_u0_u3_n143 ) , .ZN( u2_u0_u3_n168 ) );
  AND2_X1 u2_u0_u3_U80 (.A2( u2_u0_X_19 ) , .A1( u2_u0_X_20 ) , .ZN( u2_u0_u3_n104 ) );
  INV_X1 u2_u0_u3_U81 (.A( u2_u0_X_22 ) , .ZN( u2_u0_u3_n166 ) );
  INV_X1 u2_u0_u3_U82 (.A( u2_u0_X_21 ) , .ZN( u2_u0_u3_n171 ) );
  INV_X1 u2_u0_u3_U83 (.A( u2_u0_X_20 ) , .ZN( u2_u0_u3_n172 ) );
  NAND4_X1 u2_u0_u3_U84 (.ZN( u2_out0_26 ) , .A4( u2_u0_u3_n109 ) , .A3( u2_u0_u3_n110 ) , .A2( u2_u0_u3_n111 ) , .A1( u2_u0_u3_n173 ) );
  INV_X1 u2_u0_u3_U85 (.ZN( u2_u0_u3_n173 ) , .A( u2_u0_u3_n94 ) );
  OAI21_X1 u2_u0_u3_U86 (.ZN( u2_u0_u3_n111 ) , .B2( u2_u0_u3_n117 ) , .A( u2_u0_u3_n133 ) , .B1( u2_u0_u3_n176 ) );
  NAND4_X1 u2_u0_u3_U87 (.ZN( u2_out0_20 ) , .A4( u2_u0_u3_n122 ) , .A3( u2_u0_u3_n123 ) , .A1( u2_u0_u3_n175 ) , .A2( u2_u0_u3_n180 ) );
  INV_X1 u2_u0_u3_U88 (.A( u2_u0_u3_n126 ) , .ZN( u2_u0_u3_n180 ) );
  INV_X1 u2_u0_u3_U89 (.A( u2_u0_u3_n112 ) , .ZN( u2_u0_u3_n175 ) );
  OAI22_X1 u2_u0_u3_U9 (.B1( u2_u0_u3_n113 ) , .A2( u2_u0_u3_n135 ) , .A1( u2_u0_u3_n150 ) , .B2( u2_u0_u3_n164 ) , .ZN( u2_u0_u3_n98 ) );
  NAND4_X1 u2_u0_u3_U90 (.ZN( u2_out0_1 ) , .A4( u2_u0_u3_n161 ) , .A3( u2_u0_u3_n162 ) , .A2( u2_u0_u3_n163 ) , .A1( u2_u0_u3_n185 ) );
  NAND2_X1 u2_u0_u3_U91 (.ZN( u2_u0_u3_n163 ) , .A2( u2_u0_u3_n170 ) , .A1( u2_u0_u3_n176 ) );
  AOI22_X1 u2_u0_u3_U92 (.B2( u2_u0_u3_n140 ) , .B1( u2_u0_u3_n141 ) , .A2( u2_u0_u3_n142 ) , .ZN( u2_u0_u3_n162 ) , .A1( u2_u0_u3_n177 ) );
  OR4_X1 u2_u0_u3_U93 (.ZN( u2_out0_10 ) , .A4( u2_u0_u3_n136 ) , .A3( u2_u0_u3_n137 ) , .A1( u2_u0_u3_n138 ) , .A2( u2_u0_u3_n139 ) );
  OAI222_X1 u2_u0_u3_U94 (.C1( u2_u0_u3_n128 ) , .ZN( u2_u0_u3_n137 ) , .B1( u2_u0_u3_n148 ) , .A2( u2_u0_u3_n150 ) , .B2( u2_u0_u3_n154 ) , .C2( u2_u0_u3_n164 ) , .A1( u2_u0_u3_n167 ) );
  OAI221_X1 u2_u0_u3_U95 (.A( u2_u0_u3_n134 ) , .B2( u2_u0_u3_n135 ) , .ZN( u2_u0_u3_n136 ) , .C1( u2_u0_u3_n149 ) , .B1( u2_u0_u3_n151 ) , .C2( u2_u0_u3_n183 ) );
  AOI221_X1 u2_u0_u3_U96 (.A( u2_u0_u3_n131 ) , .C2( u2_u0_u3_n132 ) , .C1( u2_u0_u3_n133 ) , .ZN( u2_u0_u3_n134 ) , .B1( u2_u0_u3_n143 ) , .B2( u2_u0_u3_n177 ) );
  NAND2_X1 u2_u0_u3_U97 (.ZN( u2_u0_u3_n143 ) , .A1( u2_u0_u3_n165 ) , .A2( u2_u0_u3_n167 ) );
  NAND3_X1 u2_u0_u3_U98 (.A1( u2_u0_u3_n114 ) , .ZN( u2_u0_u3_n115 ) , .A2( u2_u0_u3_n145 ) , .A3( u2_u0_u3_n153 ) );
  NAND3_X1 u2_u0_u3_U99 (.ZN( u2_u0_u3_n129 ) , .A2( u2_u0_u3_n144 ) , .A1( u2_u0_u3_n153 ) , .A3( u2_u0_u3_n182 ) );
  OAI22_X1 u2_u0_u4_U10 (.B2( u2_u0_u4_n135 ) , .ZN( u2_u0_u4_n137 ) , .B1( u2_u0_u4_n153 ) , .A1( u2_u0_u4_n155 ) , .A2( u2_u0_u4_n171 ) );
  AND3_X1 u2_u0_u4_U11 (.A2( u2_u0_u4_n134 ) , .ZN( u2_u0_u4_n135 ) , .A3( u2_u0_u4_n145 ) , .A1( u2_u0_u4_n157 ) );
  NAND2_X1 u2_u0_u4_U12 (.ZN( u2_u0_u4_n132 ) , .A2( u2_u0_u4_n170 ) , .A1( u2_u0_u4_n173 ) );
  AOI21_X1 u2_u0_u4_U13 (.B2( u2_u0_u4_n160 ) , .B1( u2_u0_u4_n161 ) , .ZN( u2_u0_u4_n162 ) , .A( u2_u0_u4_n170 ) );
  AOI21_X1 u2_u0_u4_U14 (.ZN( u2_u0_u4_n107 ) , .B2( u2_u0_u4_n143 ) , .A( u2_u0_u4_n174 ) , .B1( u2_u0_u4_n184 ) );
  AOI21_X1 u2_u0_u4_U15 (.B2( u2_u0_u4_n158 ) , .B1( u2_u0_u4_n159 ) , .ZN( u2_u0_u4_n163 ) , .A( u2_u0_u4_n174 ) );
  AOI21_X1 u2_u0_u4_U16 (.A( u2_u0_u4_n153 ) , .B2( u2_u0_u4_n154 ) , .B1( u2_u0_u4_n155 ) , .ZN( u2_u0_u4_n165 ) );
  AOI21_X1 u2_u0_u4_U17 (.A( u2_u0_u4_n156 ) , .B2( u2_u0_u4_n157 ) , .ZN( u2_u0_u4_n164 ) , .B1( u2_u0_u4_n184 ) );
  INV_X1 u2_u0_u4_U18 (.A( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n170 ) );
  AND2_X1 u2_u0_u4_U19 (.A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n155 ) , .A1( u2_u0_u4_n160 ) );
  INV_X1 u2_u0_u4_U20 (.A( u2_u0_u4_n156 ) , .ZN( u2_u0_u4_n175 ) );
  NAND2_X1 u2_u0_u4_U21 (.A2( u2_u0_u4_n118 ) , .ZN( u2_u0_u4_n131 ) , .A1( u2_u0_u4_n147 ) );
  NAND2_X1 u2_u0_u4_U22 (.A1( u2_u0_u4_n119 ) , .A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n130 ) );
  NAND2_X1 u2_u0_u4_U23 (.ZN( u2_u0_u4_n117 ) , .A2( u2_u0_u4_n118 ) , .A1( u2_u0_u4_n148 ) );
  NAND2_X1 u2_u0_u4_U24 (.ZN( u2_u0_u4_n129 ) , .A1( u2_u0_u4_n134 ) , .A2( u2_u0_u4_n148 ) );
  AND3_X1 u2_u0_u4_U25 (.A1( u2_u0_u4_n119 ) , .A2( u2_u0_u4_n143 ) , .A3( u2_u0_u4_n154 ) , .ZN( u2_u0_u4_n161 ) );
  AND2_X1 u2_u0_u4_U26 (.A1( u2_u0_u4_n145 ) , .A2( u2_u0_u4_n147 ) , .ZN( u2_u0_u4_n159 ) );
  OR3_X1 u2_u0_u4_U27 (.A3( u2_u0_u4_n114 ) , .A2( u2_u0_u4_n115 ) , .A1( u2_u0_u4_n116 ) , .ZN( u2_u0_u4_n136 ) );
  AOI21_X1 u2_u0_u4_U28 (.A( u2_u0_u4_n113 ) , .ZN( u2_u0_u4_n116 ) , .B2( u2_u0_u4_n173 ) , .B1( u2_u0_u4_n174 ) );
  AOI21_X1 u2_u0_u4_U29 (.ZN( u2_u0_u4_n115 ) , .B2( u2_u0_u4_n145 ) , .B1( u2_u0_u4_n146 ) , .A( u2_u0_u4_n156 ) );
  NOR2_X1 u2_u0_u4_U3 (.ZN( u2_u0_u4_n121 ) , .A1( u2_u0_u4_n181 ) , .A2( u2_u0_u4_n182 ) );
  OAI22_X1 u2_u0_u4_U30 (.ZN( u2_u0_u4_n114 ) , .A2( u2_u0_u4_n121 ) , .B1( u2_u0_u4_n160 ) , .B2( u2_u0_u4_n170 ) , .A1( u2_u0_u4_n171 ) );
  INV_X1 u2_u0_u4_U31 (.A( u2_u0_u4_n158 ) , .ZN( u2_u0_u4_n182 ) );
  INV_X1 u2_u0_u4_U32 (.ZN( u2_u0_u4_n181 ) , .A( u2_u0_u4_n96 ) );
  INV_X1 u2_u0_u4_U33 (.A( u2_u0_u4_n144 ) , .ZN( u2_u0_u4_n179 ) );
  INV_X1 u2_u0_u4_U34 (.A( u2_u0_u4_n157 ) , .ZN( u2_u0_u4_n178 ) );
  NAND2_X1 u2_u0_u4_U35 (.A2( u2_u0_u4_n154 ) , .A1( u2_u0_u4_n96 ) , .ZN( u2_u0_u4_n97 ) );
  INV_X1 u2_u0_u4_U36 (.ZN( u2_u0_u4_n186 ) , .A( u2_u0_u4_n95 ) );
  OAI221_X1 u2_u0_u4_U37 (.C1( u2_u0_u4_n134 ) , .B1( u2_u0_u4_n158 ) , .B2( u2_u0_u4_n171 ) , .C2( u2_u0_u4_n173 ) , .A( u2_u0_u4_n94 ) , .ZN( u2_u0_u4_n95 ) );
  AOI222_X1 u2_u0_u4_U38 (.B2( u2_u0_u4_n132 ) , .A1( u2_u0_u4_n138 ) , .C2( u2_u0_u4_n175 ) , .A2( u2_u0_u4_n179 ) , .C1( u2_u0_u4_n181 ) , .B1( u2_u0_u4_n185 ) , .ZN( u2_u0_u4_n94 ) );
  INV_X1 u2_u0_u4_U39 (.A( u2_u0_u4_n113 ) , .ZN( u2_u0_u4_n185 ) );
  INV_X1 u2_u0_u4_U4 (.A( u2_u0_u4_n117 ) , .ZN( u2_u0_u4_n184 ) );
  INV_X1 u2_u0_u4_U40 (.A( u2_u0_u4_n143 ) , .ZN( u2_u0_u4_n183 ) );
  NOR2_X1 u2_u0_u4_U41 (.ZN( u2_u0_u4_n138 ) , .A1( u2_u0_u4_n168 ) , .A2( u2_u0_u4_n169 ) );
  NOR2_X1 u2_u0_u4_U42 (.A1( u2_u0_u4_n150 ) , .A2( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n153 ) );
  NOR2_X1 u2_u0_u4_U43 (.A2( u2_u0_u4_n128 ) , .A1( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n156 ) );
  AOI22_X1 u2_u0_u4_U44 (.B2( u2_u0_u4_n122 ) , .A1( u2_u0_u4_n123 ) , .ZN( u2_u0_u4_n124 ) , .B1( u2_u0_u4_n128 ) , .A2( u2_u0_u4_n172 ) );
  INV_X1 u2_u0_u4_U45 (.A( u2_u0_u4_n153 ) , .ZN( u2_u0_u4_n172 ) );
  NAND2_X1 u2_u0_u4_U46 (.A2( u2_u0_u4_n120 ) , .ZN( u2_u0_u4_n123 ) , .A1( u2_u0_u4_n161 ) );
  AOI22_X1 u2_u0_u4_U47 (.B2( u2_u0_u4_n132 ) , .A2( u2_u0_u4_n133 ) , .ZN( u2_u0_u4_n140 ) , .A1( u2_u0_u4_n150 ) , .B1( u2_u0_u4_n179 ) );
  NAND2_X1 u2_u0_u4_U48 (.ZN( u2_u0_u4_n133 ) , .A2( u2_u0_u4_n146 ) , .A1( u2_u0_u4_n154 ) );
  NAND2_X1 u2_u0_u4_U49 (.A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n154 ) , .A2( u2_u0_u4_n98 ) );
  NOR4_X1 u2_u0_u4_U5 (.A4( u2_u0_u4_n106 ) , .A3( u2_u0_u4_n107 ) , .A2( u2_u0_u4_n108 ) , .A1( u2_u0_u4_n109 ) , .ZN( u2_u0_u4_n110 ) );
  NAND2_X1 u2_u0_u4_U50 (.A1( u2_u0_u4_n101 ) , .ZN( u2_u0_u4_n158 ) , .A2( u2_u0_u4_n99 ) );
  AOI21_X1 u2_u0_u4_U51 (.ZN( u2_u0_u4_n127 ) , .A( u2_u0_u4_n136 ) , .B2( u2_u0_u4_n150 ) , .B1( u2_u0_u4_n180 ) );
  INV_X1 u2_u0_u4_U52 (.A( u2_u0_u4_n160 ) , .ZN( u2_u0_u4_n180 ) );
  NAND2_X1 u2_u0_u4_U53 (.A2( u2_u0_u4_n104 ) , .A1( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n146 ) );
  NAND2_X1 u2_u0_u4_U54 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n160 ) );
  NAND2_X1 u2_u0_u4_U55 (.ZN( u2_u0_u4_n134 ) , .A1( u2_u0_u4_n98 ) , .A2( u2_u0_u4_n99 ) );
  NAND2_X1 u2_u0_u4_U56 (.A1( u2_u0_u4_n103 ) , .A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n143 ) );
  NAND2_X1 u2_u0_u4_U57 (.A2( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n145 ) , .A1( u2_u0_u4_n98 ) );
  NAND2_X1 u2_u0_u4_U58 (.A1( u2_u0_u4_n100 ) , .A2( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n120 ) );
  NAND2_X1 u2_u0_u4_U59 (.A1( u2_u0_u4_n102 ) , .A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n148 ) );
  AOI21_X1 u2_u0_u4_U6 (.ZN( u2_u0_u4_n106 ) , .B2( u2_u0_u4_n146 ) , .B1( u2_u0_u4_n158 ) , .A( u2_u0_u4_n170 ) );
  NAND2_X1 u2_u0_u4_U60 (.A2( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n157 ) );
  INV_X1 u2_u0_u4_U61 (.A( u2_u0_u4_n150 ) , .ZN( u2_u0_u4_n173 ) );
  INV_X1 u2_u0_u4_U62 (.A( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n171 ) );
  NAND2_X1 u2_u0_u4_U63 (.A1( u2_u0_u4_n100 ) , .ZN( u2_u0_u4_n118 ) , .A2( u2_u0_u4_n99 ) );
  NAND2_X1 u2_u0_u4_U64 (.A2( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n144 ) );
  NAND2_X1 u2_u0_u4_U65 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n105 ) , .ZN( u2_u0_u4_n96 ) );
  INV_X1 u2_u0_u4_U66 (.A( u2_u0_u4_n128 ) , .ZN( u2_u0_u4_n174 ) );
  NAND2_X1 u2_u0_u4_U67 (.A2( u2_u0_u4_n102 ) , .ZN( u2_u0_u4_n119 ) , .A1( u2_u0_u4_n98 ) );
  NAND2_X1 u2_u0_u4_U68 (.A2( u2_u0_u4_n101 ) , .A1( u2_u0_u4_n103 ) , .ZN( u2_u0_u4_n147 ) );
  NAND2_X1 u2_u0_u4_U69 (.A2( u2_u0_u4_n104 ) , .ZN( u2_u0_u4_n113 ) , .A1( u2_u0_u4_n99 ) );
  AOI21_X1 u2_u0_u4_U7 (.ZN( u2_u0_u4_n108 ) , .B2( u2_u0_u4_n134 ) , .B1( u2_u0_u4_n155 ) , .A( u2_u0_u4_n156 ) );
  NOR2_X1 u2_u0_u4_U70 (.A2( u2_u0_X_28 ) , .ZN( u2_u0_u4_n150 ) , .A1( u2_u0_u4_n168 ) );
  NOR2_X1 u2_u0_u4_U71 (.A2( u2_u0_X_29 ) , .ZN( u2_u0_u4_n152 ) , .A1( u2_u0_u4_n169 ) );
  NOR2_X1 u2_u0_u4_U72 (.A2( u2_u0_X_30 ) , .ZN( u2_u0_u4_n105 ) , .A1( u2_u0_u4_n176 ) );
  NOR2_X1 u2_u0_u4_U73 (.A2( u2_u0_X_26 ) , .ZN( u2_u0_u4_n100 ) , .A1( u2_u0_u4_n177 ) );
  NOR2_X1 u2_u0_u4_U74 (.A2( u2_u0_X_28 ) , .A1( u2_u0_X_29 ) , .ZN( u2_u0_u4_n128 ) );
  NOR2_X1 u2_u0_u4_U75 (.A2( u2_u0_X_27 ) , .A1( u2_u0_X_30 ) , .ZN( u2_u0_u4_n102 ) );
  NOR2_X1 u2_u0_u4_U76 (.A2( u2_u0_X_25 ) , .A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n98 ) );
  AND2_X1 u2_u0_u4_U77 (.A2( u2_u0_X_25 ) , .A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n104 ) );
  AND2_X1 u2_u0_u4_U78 (.A1( u2_u0_X_30 ) , .A2( u2_u0_u4_n176 ) , .ZN( u2_u0_u4_n99 ) );
  AND2_X1 u2_u0_u4_U79 (.A1( u2_u0_X_26 ) , .ZN( u2_u0_u4_n101 ) , .A2( u2_u0_u4_n177 ) );
  AOI21_X1 u2_u0_u4_U8 (.ZN( u2_u0_u4_n109 ) , .A( u2_u0_u4_n153 ) , .B1( u2_u0_u4_n159 ) , .B2( u2_u0_u4_n184 ) );
  AND2_X1 u2_u0_u4_U80 (.A1( u2_u0_X_27 ) , .A2( u2_u0_X_30 ) , .ZN( u2_u0_u4_n103 ) );
  INV_X1 u2_u0_u4_U81 (.A( u2_u0_X_28 ) , .ZN( u2_u0_u4_n169 ) );
  INV_X1 u2_u0_u4_U82 (.A( u2_u0_X_29 ) , .ZN( u2_u0_u4_n168 ) );
  INV_X1 u2_u0_u4_U83 (.A( u2_u0_X_25 ) , .ZN( u2_u0_u4_n177 ) );
  INV_X1 u2_u0_u4_U84 (.A( u2_u0_X_27 ) , .ZN( u2_u0_u4_n176 ) );
  NAND4_X1 u2_u0_u4_U85 (.ZN( u2_out0_25 ) , .A4( u2_u0_u4_n139 ) , .A3( u2_u0_u4_n140 ) , .A2( u2_u0_u4_n141 ) , .A1( u2_u0_u4_n142 ) );
  OAI21_X1 u2_u0_u4_U86 (.A( u2_u0_u4_n128 ) , .B2( u2_u0_u4_n129 ) , .B1( u2_u0_u4_n130 ) , .ZN( u2_u0_u4_n142 ) );
  OAI21_X1 u2_u0_u4_U87 (.B2( u2_u0_u4_n131 ) , .ZN( u2_u0_u4_n141 ) , .A( u2_u0_u4_n175 ) , .B1( u2_u0_u4_n183 ) );
  NAND4_X1 u2_u0_u4_U88 (.ZN( u2_out0_14 ) , .A4( u2_u0_u4_n124 ) , .A3( u2_u0_u4_n125 ) , .A2( u2_u0_u4_n126 ) , .A1( u2_u0_u4_n127 ) );
  AOI22_X1 u2_u0_u4_U89 (.B2( u2_u0_u4_n117 ) , .ZN( u2_u0_u4_n126 ) , .A1( u2_u0_u4_n129 ) , .B1( u2_u0_u4_n152 ) , .A2( u2_u0_u4_n175 ) );
  AOI211_X1 u2_u0_u4_U9 (.B( u2_u0_u4_n136 ) , .A( u2_u0_u4_n137 ) , .C2( u2_u0_u4_n138 ) , .ZN( u2_u0_u4_n139 ) , .C1( u2_u0_u4_n182 ) );
  AOI22_X1 u2_u0_u4_U90 (.ZN( u2_u0_u4_n125 ) , .B2( u2_u0_u4_n131 ) , .A2( u2_u0_u4_n132 ) , .B1( u2_u0_u4_n138 ) , .A1( u2_u0_u4_n178 ) );
  NAND4_X1 u2_u0_u4_U91 (.ZN( u2_out0_8 ) , .A4( u2_u0_u4_n110 ) , .A3( u2_u0_u4_n111 ) , .A2( u2_u0_u4_n112 ) , .A1( u2_u0_u4_n186 ) );
  NAND2_X1 u2_u0_u4_U92 (.ZN( u2_u0_u4_n112 ) , .A2( u2_u0_u4_n130 ) , .A1( u2_u0_u4_n150 ) );
  AOI22_X1 u2_u0_u4_U93 (.ZN( u2_u0_u4_n111 ) , .B2( u2_u0_u4_n132 ) , .A1( u2_u0_u4_n152 ) , .B1( u2_u0_u4_n178 ) , .A2( u2_u0_u4_n97 ) );
  AOI22_X1 u2_u0_u4_U94 (.B2( u2_u0_u4_n149 ) , .B1( u2_u0_u4_n150 ) , .A2( u2_u0_u4_n151 ) , .A1( u2_u0_u4_n152 ) , .ZN( u2_u0_u4_n167 ) );
  NOR4_X1 u2_u0_u4_U95 (.A4( u2_u0_u4_n162 ) , .A3( u2_u0_u4_n163 ) , .A2( u2_u0_u4_n164 ) , .A1( u2_u0_u4_n165 ) , .ZN( u2_u0_u4_n166 ) );
  NAND3_X1 u2_u0_u4_U96 (.ZN( u2_out0_3 ) , .A3( u2_u0_u4_n166 ) , .A1( u2_u0_u4_n167 ) , .A2( u2_u0_u4_n186 ) );
  NAND3_X1 u2_u0_u4_U97 (.A3( u2_u0_u4_n146 ) , .A2( u2_u0_u4_n147 ) , .A1( u2_u0_u4_n148 ) , .ZN( u2_u0_u4_n149 ) );
  NAND3_X1 u2_u0_u4_U98 (.A3( u2_u0_u4_n143 ) , .A2( u2_u0_u4_n144 ) , .A1( u2_u0_u4_n145 ) , .ZN( u2_u0_u4_n151 ) );
  NAND3_X1 u2_u0_u4_U99 (.A3( u2_u0_u4_n121 ) , .ZN( u2_u0_u4_n122 ) , .A2( u2_u0_u4_n144 ) , .A1( u2_u0_u4_n154 ) );
  INV_X1 u2_u0_u5_U10 (.A( u2_u0_u5_n121 ) , .ZN( u2_u0_u5_n177 ) );
  NOR3_X1 u2_u0_u5_U100 (.A3( u2_u0_u5_n141 ) , .A1( u2_u0_u5_n142 ) , .ZN( u2_u0_u5_n143 ) , .A2( u2_u0_u5_n191 ) );
  NAND4_X1 u2_u0_u5_U101 (.ZN( u2_out0_4 ) , .A4( u2_u0_u5_n112 ) , .A2( u2_u0_u5_n113 ) , .A1( u2_u0_u5_n114 ) , .A3( u2_u0_u5_n195 ) );
  AOI211_X1 u2_u0_u5_U102 (.A( u2_u0_u5_n110 ) , .C1( u2_u0_u5_n111 ) , .ZN( u2_u0_u5_n112 ) , .B( u2_u0_u5_n118 ) , .C2( u2_u0_u5_n177 ) );
  AOI222_X1 u2_u0_u5_U103 (.ZN( u2_u0_u5_n113 ) , .A1( u2_u0_u5_n131 ) , .C1( u2_u0_u5_n148 ) , .B2( u2_u0_u5_n174 ) , .C2( u2_u0_u5_n178 ) , .A2( u2_u0_u5_n179 ) , .B1( u2_u0_u5_n99 ) );
  NAND3_X1 u2_u0_u5_U104 (.A2( u2_u0_u5_n154 ) , .A3( u2_u0_u5_n158 ) , .A1( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n99 ) );
  NOR2_X1 u2_u0_u5_U11 (.ZN( u2_u0_u5_n160 ) , .A2( u2_u0_u5_n173 ) , .A1( u2_u0_u5_n177 ) );
  INV_X1 u2_u0_u5_U12 (.A( u2_u0_u5_n150 ) , .ZN( u2_u0_u5_n174 ) );
  AOI21_X1 u2_u0_u5_U13 (.A( u2_u0_u5_n160 ) , .B2( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n162 ) , .B1( u2_u0_u5_n192 ) );
  INV_X1 u2_u0_u5_U14 (.A( u2_u0_u5_n159 ) , .ZN( u2_u0_u5_n192 ) );
  AOI21_X1 u2_u0_u5_U15 (.A( u2_u0_u5_n156 ) , .B2( u2_u0_u5_n157 ) , .B1( u2_u0_u5_n158 ) , .ZN( u2_u0_u5_n163 ) );
  AOI21_X1 u2_u0_u5_U16 (.B2( u2_u0_u5_n139 ) , .B1( u2_u0_u5_n140 ) , .ZN( u2_u0_u5_n141 ) , .A( u2_u0_u5_n150 ) );
  OAI21_X1 u2_u0_u5_U17 (.A( u2_u0_u5_n133 ) , .B2( u2_u0_u5_n134 ) , .B1( u2_u0_u5_n135 ) , .ZN( u2_u0_u5_n142 ) );
  OAI21_X1 u2_u0_u5_U18 (.ZN( u2_u0_u5_n133 ) , .B2( u2_u0_u5_n147 ) , .A( u2_u0_u5_n173 ) , .B1( u2_u0_u5_n188 ) );
  NAND2_X1 u2_u0_u5_U19 (.A2( u2_u0_u5_n119 ) , .A1( u2_u0_u5_n123 ) , .ZN( u2_u0_u5_n137 ) );
  INV_X1 u2_u0_u5_U20 (.A( u2_u0_u5_n155 ) , .ZN( u2_u0_u5_n194 ) );
  NAND2_X1 u2_u0_u5_U21 (.A1( u2_u0_u5_n121 ) , .ZN( u2_u0_u5_n132 ) , .A2( u2_u0_u5_n172 ) );
  NAND2_X1 u2_u0_u5_U22 (.A2( u2_u0_u5_n122 ) , .ZN( u2_u0_u5_n136 ) , .A1( u2_u0_u5_n154 ) );
  NAND2_X1 u2_u0_u5_U23 (.A2( u2_u0_u5_n119 ) , .A1( u2_u0_u5_n120 ) , .ZN( u2_u0_u5_n159 ) );
  INV_X1 u2_u0_u5_U24 (.A( u2_u0_u5_n156 ) , .ZN( u2_u0_u5_n175 ) );
  INV_X1 u2_u0_u5_U25 (.A( u2_u0_u5_n158 ) , .ZN( u2_u0_u5_n188 ) );
  INV_X1 u2_u0_u5_U26 (.A( u2_u0_u5_n152 ) , .ZN( u2_u0_u5_n179 ) );
  INV_X1 u2_u0_u5_U27 (.A( u2_u0_u5_n140 ) , .ZN( u2_u0_u5_n182 ) );
  INV_X1 u2_u0_u5_U28 (.A( u2_u0_u5_n151 ) , .ZN( u2_u0_u5_n183 ) );
  INV_X1 u2_u0_u5_U29 (.A( u2_u0_u5_n123 ) , .ZN( u2_u0_u5_n185 ) );
  NOR2_X1 u2_u0_u5_U3 (.ZN( u2_u0_u5_n134 ) , .A1( u2_u0_u5_n183 ) , .A2( u2_u0_u5_n190 ) );
  INV_X1 u2_u0_u5_U30 (.A( u2_u0_u5_n161 ) , .ZN( u2_u0_u5_n184 ) );
  INV_X1 u2_u0_u5_U31 (.A( u2_u0_u5_n139 ) , .ZN( u2_u0_u5_n189 ) );
  INV_X1 u2_u0_u5_U32 (.A( u2_u0_u5_n157 ) , .ZN( u2_u0_u5_n190 ) );
  INV_X1 u2_u0_u5_U33 (.A( u2_u0_u5_n120 ) , .ZN( u2_u0_u5_n193 ) );
  NAND2_X1 u2_u0_u5_U34 (.ZN( u2_u0_u5_n111 ) , .A1( u2_u0_u5_n140 ) , .A2( u2_u0_u5_n155 ) );
  NOR2_X1 u2_u0_u5_U35 (.ZN( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n170 ) , .A2( u2_u0_u5_n180 ) );
  INV_X1 u2_u0_u5_U36 (.A( u2_u0_u5_n117 ) , .ZN( u2_u0_u5_n196 ) );
  OAI221_X1 u2_u0_u5_U37 (.A( u2_u0_u5_n116 ) , .ZN( u2_u0_u5_n117 ) , .B2( u2_u0_u5_n119 ) , .C1( u2_u0_u5_n153 ) , .C2( u2_u0_u5_n158 ) , .B1( u2_u0_u5_n172 ) );
  AOI222_X1 u2_u0_u5_U38 (.ZN( u2_u0_u5_n116 ) , .B2( u2_u0_u5_n145 ) , .C1( u2_u0_u5_n148 ) , .A2( u2_u0_u5_n174 ) , .C2( u2_u0_u5_n177 ) , .B1( u2_u0_u5_n187 ) , .A1( u2_u0_u5_n193 ) );
  INV_X1 u2_u0_u5_U39 (.A( u2_u0_u5_n115 ) , .ZN( u2_u0_u5_n187 ) );
  INV_X1 u2_u0_u5_U4 (.A( u2_u0_u5_n138 ) , .ZN( u2_u0_u5_n191 ) );
  AOI22_X1 u2_u0_u5_U40 (.B2( u2_u0_u5_n131 ) , .A2( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n169 ) , .B1( u2_u0_u5_n174 ) , .A1( u2_u0_u5_n185 ) );
  NOR2_X1 u2_u0_u5_U41 (.A1( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n150 ) , .A2( u2_u0_u5_n173 ) );
  AOI21_X1 u2_u0_u5_U42 (.A( u2_u0_u5_n118 ) , .B2( u2_u0_u5_n145 ) , .ZN( u2_u0_u5_n168 ) , .B1( u2_u0_u5_n186 ) );
  INV_X1 u2_u0_u5_U43 (.A( u2_u0_u5_n122 ) , .ZN( u2_u0_u5_n186 ) );
  NOR2_X1 u2_u0_u5_U44 (.A1( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n152 ) , .A2( u2_u0_u5_n176 ) );
  NOR2_X1 u2_u0_u5_U45 (.A1( u2_u0_u5_n115 ) , .ZN( u2_u0_u5_n118 ) , .A2( u2_u0_u5_n153 ) );
  NOR2_X1 u2_u0_u5_U46 (.A2( u2_u0_u5_n145 ) , .ZN( u2_u0_u5_n156 ) , .A1( u2_u0_u5_n174 ) );
  NOR2_X1 u2_u0_u5_U47 (.ZN( u2_u0_u5_n121 ) , .A2( u2_u0_u5_n145 ) , .A1( u2_u0_u5_n176 ) );
  AOI22_X1 u2_u0_u5_U48 (.ZN( u2_u0_u5_n114 ) , .A2( u2_u0_u5_n137 ) , .A1( u2_u0_u5_n145 ) , .B2( u2_u0_u5_n175 ) , .B1( u2_u0_u5_n193 ) );
  OAI211_X1 u2_u0_u5_U49 (.B( u2_u0_u5_n124 ) , .A( u2_u0_u5_n125 ) , .C2( u2_u0_u5_n126 ) , .C1( u2_u0_u5_n127 ) , .ZN( u2_u0_u5_n128 ) );
  OAI21_X1 u2_u0_u5_U5 (.B2( u2_u0_u5_n136 ) , .B1( u2_u0_u5_n137 ) , .ZN( u2_u0_u5_n138 ) , .A( u2_u0_u5_n177 ) );
  NOR3_X1 u2_u0_u5_U50 (.ZN( u2_u0_u5_n127 ) , .A1( u2_u0_u5_n136 ) , .A3( u2_u0_u5_n148 ) , .A2( u2_u0_u5_n182 ) );
  OAI21_X1 u2_u0_u5_U51 (.ZN( u2_u0_u5_n124 ) , .A( u2_u0_u5_n177 ) , .B2( u2_u0_u5_n183 ) , .B1( u2_u0_u5_n189 ) );
  OAI21_X1 u2_u0_u5_U52 (.ZN( u2_u0_u5_n125 ) , .A( u2_u0_u5_n174 ) , .B2( u2_u0_u5_n185 ) , .B1( u2_u0_u5_n190 ) );
  AOI21_X1 u2_u0_u5_U53 (.A( u2_u0_u5_n153 ) , .B2( u2_u0_u5_n154 ) , .B1( u2_u0_u5_n155 ) , .ZN( u2_u0_u5_n164 ) );
  AOI21_X1 u2_u0_u5_U54 (.ZN( u2_u0_u5_n110 ) , .B1( u2_u0_u5_n122 ) , .B2( u2_u0_u5_n139 ) , .A( u2_u0_u5_n153 ) );
  INV_X1 u2_u0_u5_U55 (.A( u2_u0_u5_n153 ) , .ZN( u2_u0_u5_n176 ) );
  INV_X1 u2_u0_u5_U56 (.A( u2_u0_u5_n126 ) , .ZN( u2_u0_u5_n173 ) );
  AND2_X1 u2_u0_u5_U57 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n147 ) );
  AND2_X1 u2_u0_u5_U58 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n148 ) );
  NAND2_X1 u2_u0_u5_U59 (.A1( u2_u0_u5_n105 ) , .A2( u2_u0_u5_n106 ) , .ZN( u2_u0_u5_n158 ) );
  INV_X1 u2_u0_u5_U6 (.A( u2_u0_u5_n135 ) , .ZN( u2_u0_u5_n178 ) );
  NAND2_X1 u2_u0_u5_U60 (.A2( u2_u0_u5_n108 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n139 ) );
  NAND2_X1 u2_u0_u5_U61 (.A1( u2_u0_u5_n106 ) , .A2( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n119 ) );
  NAND2_X1 u2_u0_u5_U62 (.A2( u2_u0_u5_n103 ) , .A1( u2_u0_u5_n105 ) , .ZN( u2_u0_u5_n140 ) );
  NAND2_X1 u2_u0_u5_U63 (.A2( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n105 ) , .ZN( u2_u0_u5_n155 ) );
  NAND2_X1 u2_u0_u5_U64 (.A2( u2_u0_u5_n106 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n122 ) );
  NAND2_X1 u2_u0_u5_U65 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n106 ) , .ZN( u2_u0_u5_n115 ) );
  NAND2_X1 u2_u0_u5_U66 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n103 ) , .ZN( u2_u0_u5_n161 ) );
  NAND2_X1 u2_u0_u5_U67 (.A1( u2_u0_u5_n105 ) , .A2( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n154 ) );
  INV_X1 u2_u0_u5_U68 (.A( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n172 ) );
  NAND2_X1 u2_u0_u5_U69 (.A1( u2_u0_u5_n103 ) , .A2( u2_u0_u5_n108 ) , .ZN( u2_u0_u5_n123 ) );
  OAI22_X1 u2_u0_u5_U7 (.B2( u2_u0_u5_n149 ) , .B1( u2_u0_u5_n150 ) , .A2( u2_u0_u5_n151 ) , .A1( u2_u0_u5_n152 ) , .ZN( u2_u0_u5_n165 ) );
  NAND2_X1 u2_u0_u5_U70 (.A2( u2_u0_u5_n103 ) , .A1( u2_u0_u5_n107 ) , .ZN( u2_u0_u5_n151 ) );
  NAND2_X1 u2_u0_u5_U71 (.A2( u2_u0_u5_n107 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n120 ) );
  NAND2_X1 u2_u0_u5_U72 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n109 ) , .ZN( u2_u0_u5_n157 ) );
  AND2_X1 u2_u0_u5_U73 (.A2( u2_u0_u5_n100 ) , .A1( u2_u0_u5_n104 ) , .ZN( u2_u0_u5_n131 ) );
  INV_X1 u2_u0_u5_U74 (.A( u2_u0_u5_n102 ) , .ZN( u2_u0_u5_n195 ) );
  OAI221_X1 u2_u0_u5_U75 (.A( u2_u0_u5_n101 ) , .ZN( u2_u0_u5_n102 ) , .C2( u2_u0_u5_n115 ) , .C1( u2_u0_u5_n126 ) , .B1( u2_u0_u5_n134 ) , .B2( u2_u0_u5_n160 ) );
  OAI21_X1 u2_u0_u5_U76 (.ZN( u2_u0_u5_n101 ) , .B1( u2_u0_u5_n137 ) , .A( u2_u0_u5_n146 ) , .B2( u2_u0_u5_n147 ) );
  NOR2_X1 u2_u0_u5_U77 (.A2( u2_u0_X_34 ) , .A1( u2_u0_X_35 ) , .ZN( u2_u0_u5_n145 ) );
  NOR2_X1 u2_u0_u5_U78 (.A2( u2_u0_X_34 ) , .ZN( u2_u0_u5_n146 ) , .A1( u2_u0_u5_n171 ) );
  NOR2_X1 u2_u0_u5_U79 (.A2( u2_u0_X_31 ) , .A1( u2_u0_X_32 ) , .ZN( u2_u0_u5_n103 ) );
  NOR3_X1 u2_u0_u5_U8 (.A2( u2_u0_u5_n147 ) , .A1( u2_u0_u5_n148 ) , .ZN( u2_u0_u5_n149 ) , .A3( u2_u0_u5_n194 ) );
  NOR2_X1 u2_u0_u5_U80 (.A2( u2_u0_X_36 ) , .ZN( u2_u0_u5_n105 ) , .A1( u2_u0_u5_n180 ) );
  NOR2_X1 u2_u0_u5_U81 (.A2( u2_u0_X_33 ) , .ZN( u2_u0_u5_n108 ) , .A1( u2_u0_u5_n170 ) );
  NOR2_X1 u2_u0_u5_U82 (.A2( u2_u0_X_33 ) , .A1( u2_u0_X_36 ) , .ZN( u2_u0_u5_n107 ) );
  NOR2_X1 u2_u0_u5_U83 (.A2( u2_u0_X_31 ) , .ZN( u2_u0_u5_n104 ) , .A1( u2_u0_u5_n181 ) );
  NAND2_X1 u2_u0_u5_U84 (.A2( u2_u0_X_34 ) , .A1( u2_u0_X_35 ) , .ZN( u2_u0_u5_n153 ) );
  NAND2_X1 u2_u0_u5_U85 (.A1( u2_u0_X_34 ) , .ZN( u2_u0_u5_n126 ) , .A2( u2_u0_u5_n171 ) );
  AND2_X1 u2_u0_u5_U86 (.A1( u2_u0_X_31 ) , .A2( u2_u0_X_32 ) , .ZN( u2_u0_u5_n106 ) );
  AND2_X1 u2_u0_u5_U87 (.A1( u2_u0_X_31 ) , .ZN( u2_u0_u5_n109 ) , .A2( u2_u0_u5_n181 ) );
  INV_X1 u2_u0_u5_U88 (.A( u2_u0_X_33 ) , .ZN( u2_u0_u5_n180 ) );
  INV_X1 u2_u0_u5_U89 (.A( u2_u0_X_35 ) , .ZN( u2_u0_u5_n171 ) );
  NOR2_X1 u2_u0_u5_U9 (.ZN( u2_u0_u5_n135 ) , .A1( u2_u0_u5_n173 ) , .A2( u2_u0_u5_n176 ) );
  INV_X1 u2_u0_u5_U90 (.A( u2_u0_X_36 ) , .ZN( u2_u0_u5_n170 ) );
  INV_X1 u2_u0_u5_U91 (.A( u2_u0_X_32 ) , .ZN( u2_u0_u5_n181 ) );
  NAND4_X1 u2_u0_u5_U92 (.ZN( u2_out0_29 ) , .A4( u2_u0_u5_n129 ) , .A3( u2_u0_u5_n130 ) , .A2( u2_u0_u5_n168 ) , .A1( u2_u0_u5_n196 ) );
  AOI221_X1 u2_u0_u5_U93 (.A( u2_u0_u5_n128 ) , .ZN( u2_u0_u5_n129 ) , .C2( u2_u0_u5_n132 ) , .B2( u2_u0_u5_n159 ) , .B1( u2_u0_u5_n176 ) , .C1( u2_u0_u5_n184 ) );
  AOI222_X1 u2_u0_u5_U94 (.ZN( u2_u0_u5_n130 ) , .A2( u2_u0_u5_n146 ) , .B1( u2_u0_u5_n147 ) , .C2( u2_u0_u5_n175 ) , .B2( u2_u0_u5_n179 ) , .A1( u2_u0_u5_n188 ) , .C1( u2_u0_u5_n194 ) );
  NAND4_X1 u2_u0_u5_U95 (.ZN( u2_out0_19 ) , .A4( u2_u0_u5_n166 ) , .A3( u2_u0_u5_n167 ) , .A2( u2_u0_u5_n168 ) , .A1( u2_u0_u5_n169 ) );
  AOI22_X1 u2_u0_u5_U96 (.B2( u2_u0_u5_n145 ) , .A2( u2_u0_u5_n146 ) , .ZN( u2_u0_u5_n167 ) , .B1( u2_u0_u5_n182 ) , .A1( u2_u0_u5_n189 ) );
  NOR4_X1 u2_u0_u5_U97 (.A4( u2_u0_u5_n162 ) , .A3( u2_u0_u5_n163 ) , .A2( u2_u0_u5_n164 ) , .A1( u2_u0_u5_n165 ) , .ZN( u2_u0_u5_n166 ) );
  NAND4_X1 u2_u0_u5_U98 (.ZN( u2_out0_11 ) , .A4( u2_u0_u5_n143 ) , .A3( u2_u0_u5_n144 ) , .A2( u2_u0_u5_n169 ) , .A1( u2_u0_u5_n196 ) );
  AOI22_X1 u2_u0_u5_U99 (.A2( u2_u0_u5_n132 ) , .ZN( u2_u0_u5_n144 ) , .B2( u2_u0_u5_n145 ) , .B1( u2_u0_u5_n184 ) , .A1( u2_u0_u5_n194 ) );
  AOI22_X1 u2_u0_u6_U10 (.A2( u2_u0_u6_n151 ) , .B2( u2_u0_u6_n161 ) , .A1( u2_u0_u6_n167 ) , .B1( u2_u0_u6_n170 ) , .ZN( u2_u0_u6_n89 ) );
  AOI21_X1 u2_u0_u6_U11 (.B1( u2_u0_u6_n107 ) , .B2( u2_u0_u6_n132 ) , .A( u2_u0_u6_n158 ) , .ZN( u2_u0_u6_n88 ) );
  AOI21_X1 u2_u0_u6_U12 (.B2( u2_u0_u6_n147 ) , .B1( u2_u0_u6_n148 ) , .ZN( u2_u0_u6_n149 ) , .A( u2_u0_u6_n158 ) );
  AOI21_X1 u2_u0_u6_U13 (.ZN( u2_u0_u6_n106 ) , .A( u2_u0_u6_n142 ) , .B2( u2_u0_u6_n159 ) , .B1( u2_u0_u6_n164 ) );
  INV_X1 u2_u0_u6_U14 (.A( u2_u0_u6_n155 ) , .ZN( u2_u0_u6_n161 ) );
  INV_X1 u2_u0_u6_U15 (.A( u2_u0_u6_n128 ) , .ZN( u2_u0_u6_n164 ) );
  NAND2_X1 u2_u0_u6_U16 (.ZN( u2_u0_u6_n110 ) , .A1( u2_u0_u6_n122 ) , .A2( u2_u0_u6_n129 ) );
  NAND2_X1 u2_u0_u6_U17 (.ZN( u2_u0_u6_n124 ) , .A2( u2_u0_u6_n146 ) , .A1( u2_u0_u6_n148 ) );
  INV_X1 u2_u0_u6_U18 (.A( u2_u0_u6_n132 ) , .ZN( u2_u0_u6_n171 ) );
  AND2_X1 u2_u0_u6_U19 (.A1( u2_u0_u6_n100 ) , .ZN( u2_u0_u6_n130 ) , .A2( u2_u0_u6_n147 ) );
  INV_X1 u2_u0_u6_U20 (.A( u2_u0_u6_n127 ) , .ZN( u2_u0_u6_n173 ) );
  INV_X1 u2_u0_u6_U21 (.A( u2_u0_u6_n121 ) , .ZN( u2_u0_u6_n167 ) );
  INV_X1 u2_u0_u6_U22 (.A( u2_u0_u6_n100 ) , .ZN( u2_u0_u6_n169 ) );
  INV_X1 u2_u0_u6_U23 (.A( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n170 ) );
  INV_X1 u2_u0_u6_U24 (.A( u2_u0_u6_n113 ) , .ZN( u2_u0_u6_n168 ) );
  AND2_X1 u2_u0_u6_U25 (.A1( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n119 ) , .ZN( u2_u0_u6_n133 ) );
  AND2_X1 u2_u0_u6_U26 (.A2( u2_u0_u6_n121 ) , .A1( u2_u0_u6_n122 ) , .ZN( u2_u0_u6_n131 ) );
  AND3_X1 u2_u0_u6_U27 (.ZN( u2_u0_u6_n120 ) , .A2( u2_u0_u6_n127 ) , .A1( u2_u0_u6_n132 ) , .A3( u2_u0_u6_n145 ) );
  INV_X1 u2_u0_u6_U28 (.A( u2_u0_u6_n146 ) , .ZN( u2_u0_u6_n163 ) );
  AOI222_X1 u2_u0_u6_U29 (.ZN( u2_u0_u6_n114 ) , .A1( u2_u0_u6_n118 ) , .A2( u2_u0_u6_n126 ) , .B2( u2_u0_u6_n151 ) , .C2( u2_u0_u6_n159 ) , .C1( u2_u0_u6_n168 ) , .B1( u2_u0_u6_n169 ) );
  INV_X1 u2_u0_u6_U3 (.A( u2_u0_u6_n110 ) , .ZN( u2_u0_u6_n166 ) );
  NOR2_X1 u2_u0_u6_U30 (.A1( u2_u0_u6_n162 ) , .A2( u2_u0_u6_n165 ) , .ZN( u2_u0_u6_n98 ) );
  AOI211_X1 u2_u0_u6_U31 (.B( u2_u0_u6_n134 ) , .A( u2_u0_u6_n135 ) , .C1( u2_u0_u6_n136 ) , .ZN( u2_u0_u6_n137 ) , .C2( u2_u0_u6_n151 ) );
  AOI21_X1 u2_u0_u6_U32 (.B2( u2_u0_u6_n132 ) , .B1( u2_u0_u6_n133 ) , .ZN( u2_u0_u6_n134 ) , .A( u2_u0_u6_n158 ) );
  NAND4_X1 u2_u0_u6_U33 (.A4( u2_u0_u6_n127 ) , .A3( u2_u0_u6_n128 ) , .A2( u2_u0_u6_n129 ) , .A1( u2_u0_u6_n130 ) , .ZN( u2_u0_u6_n136 ) );
  AOI21_X1 u2_u0_u6_U34 (.B1( u2_u0_u6_n131 ) , .ZN( u2_u0_u6_n135 ) , .A( u2_u0_u6_n144 ) , .B2( u2_u0_u6_n146 ) );
  NAND2_X1 u2_u0_u6_U35 (.A1( u2_u0_u6_n144 ) , .ZN( u2_u0_u6_n151 ) , .A2( u2_u0_u6_n158 ) );
  NAND2_X1 u2_u0_u6_U36 (.ZN( u2_u0_u6_n132 ) , .A1( u2_u0_u6_n91 ) , .A2( u2_u0_u6_n97 ) );
  AOI22_X1 u2_u0_u6_U37 (.B2( u2_u0_u6_n110 ) , .B1( u2_u0_u6_n111 ) , .A1( u2_u0_u6_n112 ) , .ZN( u2_u0_u6_n115 ) , .A2( u2_u0_u6_n161 ) );
  NAND4_X1 u2_u0_u6_U38 (.A3( u2_u0_u6_n109 ) , .ZN( u2_u0_u6_n112 ) , .A4( u2_u0_u6_n132 ) , .A2( u2_u0_u6_n147 ) , .A1( u2_u0_u6_n166 ) );
  NOR2_X1 u2_u0_u6_U39 (.ZN( u2_u0_u6_n109 ) , .A1( u2_u0_u6_n170 ) , .A2( u2_u0_u6_n173 ) );
  INV_X1 u2_u0_u6_U4 (.A( u2_u0_u6_n142 ) , .ZN( u2_u0_u6_n174 ) );
  NOR2_X1 u2_u0_u6_U40 (.A2( u2_u0_u6_n126 ) , .ZN( u2_u0_u6_n155 ) , .A1( u2_u0_u6_n160 ) );
  NAND2_X1 u2_u0_u6_U41 (.ZN( u2_u0_u6_n146 ) , .A2( u2_u0_u6_n94 ) , .A1( u2_u0_u6_n99 ) );
  AOI21_X1 u2_u0_u6_U42 (.A( u2_u0_u6_n144 ) , .B2( u2_u0_u6_n145 ) , .B1( u2_u0_u6_n146 ) , .ZN( u2_u0_u6_n150 ) );
  INV_X1 u2_u0_u6_U43 (.A( u2_u0_u6_n111 ) , .ZN( u2_u0_u6_n158 ) );
  NAND2_X1 u2_u0_u6_U44 (.ZN( u2_u0_u6_n127 ) , .A1( u2_u0_u6_n91 ) , .A2( u2_u0_u6_n92 ) );
  NAND2_X1 u2_u0_u6_U45 (.ZN( u2_u0_u6_n129 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n96 ) );
  INV_X1 u2_u0_u6_U46 (.A( u2_u0_u6_n144 ) , .ZN( u2_u0_u6_n159 ) );
  NAND2_X1 u2_u0_u6_U47 (.ZN( u2_u0_u6_n145 ) , .A2( u2_u0_u6_n97 ) , .A1( u2_u0_u6_n98 ) );
  NAND2_X1 u2_u0_u6_U48 (.ZN( u2_u0_u6_n148 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n94 ) );
  NAND2_X1 u2_u0_u6_U49 (.ZN( u2_u0_u6_n108 ) , .A2( u2_u0_u6_n139 ) , .A1( u2_u0_u6_n144 ) );
  NAND2_X1 u2_u0_u6_U5 (.A2( u2_u0_u6_n143 ) , .ZN( u2_u0_u6_n152 ) , .A1( u2_u0_u6_n166 ) );
  NAND2_X1 u2_u0_u6_U50 (.ZN( u2_u0_u6_n121 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n97 ) );
  NAND2_X1 u2_u0_u6_U51 (.ZN( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n95 ) );
  AND2_X1 u2_u0_u6_U52 (.ZN( u2_u0_u6_n118 ) , .A2( u2_u0_u6_n91 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U53 (.ZN( u2_u0_u6_n147 ) , .A2( u2_u0_u6_n98 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U54 (.ZN( u2_u0_u6_n128 ) , .A1( u2_u0_u6_n94 ) , .A2( u2_u0_u6_n96 ) );
  NAND2_X1 u2_u0_u6_U55 (.ZN( u2_u0_u6_n119 ) , .A2( u2_u0_u6_n95 ) , .A1( u2_u0_u6_n99 ) );
  NAND2_X1 u2_u0_u6_U56 (.ZN( u2_u0_u6_n123 ) , .A2( u2_u0_u6_n91 ) , .A1( u2_u0_u6_n96 ) );
  NAND2_X1 u2_u0_u6_U57 (.ZN( u2_u0_u6_n100 ) , .A2( u2_u0_u6_n92 ) , .A1( u2_u0_u6_n98 ) );
  NAND2_X1 u2_u0_u6_U58 (.ZN( u2_u0_u6_n122 ) , .A1( u2_u0_u6_n94 ) , .A2( u2_u0_u6_n97 ) );
  INV_X1 u2_u0_u6_U59 (.A( u2_u0_u6_n139 ) , .ZN( u2_u0_u6_n160 ) );
  AOI22_X1 u2_u0_u6_U6 (.B2( u2_u0_u6_n101 ) , .A1( u2_u0_u6_n102 ) , .ZN( u2_u0_u6_n103 ) , .B1( u2_u0_u6_n160 ) , .A2( u2_u0_u6_n161 ) );
  NAND2_X1 u2_u0_u6_U60 (.ZN( u2_u0_u6_n113 ) , .A1( u2_u0_u6_n96 ) , .A2( u2_u0_u6_n98 ) );
  NOR2_X1 u2_u0_u6_U61 (.A2( u2_u0_X_40 ) , .A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n126 ) );
  NOR2_X1 u2_u0_u6_U62 (.A2( u2_u0_X_39 ) , .A1( u2_u0_X_42 ) , .ZN( u2_u0_u6_n92 ) );
  NOR2_X1 u2_u0_u6_U63 (.A2( u2_u0_X_39 ) , .A1( u2_u0_u6_n156 ) , .ZN( u2_u0_u6_n97 ) );
  NOR2_X1 u2_u0_u6_U64 (.A2( u2_u0_X_38 ) , .A1( u2_u0_u6_n165 ) , .ZN( u2_u0_u6_n95 ) );
  NOR2_X1 u2_u0_u6_U65 (.A2( u2_u0_X_41 ) , .ZN( u2_u0_u6_n111 ) , .A1( u2_u0_u6_n157 ) );
  NOR2_X1 u2_u0_u6_U66 (.A2( u2_u0_X_37 ) , .A1( u2_u0_u6_n162 ) , .ZN( u2_u0_u6_n94 ) );
  NOR2_X1 u2_u0_u6_U67 (.A2( u2_u0_X_37 ) , .A1( u2_u0_X_38 ) , .ZN( u2_u0_u6_n91 ) );
  NAND2_X1 u2_u0_u6_U68 (.A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n144 ) , .A2( u2_u0_u6_n157 ) );
  NAND2_X1 u2_u0_u6_U69 (.A2( u2_u0_X_40 ) , .A1( u2_u0_X_41 ) , .ZN( u2_u0_u6_n139 ) );
  NOR2_X1 u2_u0_u6_U7 (.A1( u2_u0_u6_n118 ) , .ZN( u2_u0_u6_n143 ) , .A2( u2_u0_u6_n168 ) );
  AND2_X1 u2_u0_u6_U70 (.A1( u2_u0_X_39 ) , .A2( u2_u0_u6_n156 ) , .ZN( u2_u0_u6_n96 ) );
  AND2_X1 u2_u0_u6_U71 (.A1( u2_u0_X_39 ) , .A2( u2_u0_X_42 ) , .ZN( u2_u0_u6_n99 ) );
  INV_X1 u2_u0_u6_U72 (.A( u2_u0_X_40 ) , .ZN( u2_u0_u6_n157 ) );
  INV_X1 u2_u0_u6_U73 (.A( u2_u0_X_37 ) , .ZN( u2_u0_u6_n165 ) );
  INV_X1 u2_u0_u6_U74 (.A( u2_u0_X_38 ) , .ZN( u2_u0_u6_n162 ) );
  INV_X1 u2_u0_u6_U75 (.A( u2_u0_X_42 ) , .ZN( u2_u0_u6_n156 ) );
  NAND4_X1 u2_u0_u6_U76 (.ZN( u2_out0_32 ) , .A4( u2_u0_u6_n103 ) , .A3( u2_u0_u6_n104 ) , .A2( u2_u0_u6_n105 ) , .A1( u2_u0_u6_n106 ) );
  AOI22_X1 u2_u0_u6_U77 (.ZN( u2_u0_u6_n105 ) , .A2( u2_u0_u6_n108 ) , .A1( u2_u0_u6_n118 ) , .B2( u2_u0_u6_n126 ) , .B1( u2_u0_u6_n171 ) );
  AOI22_X1 u2_u0_u6_U78 (.ZN( u2_u0_u6_n104 ) , .A1( u2_u0_u6_n111 ) , .B1( u2_u0_u6_n124 ) , .B2( u2_u0_u6_n151 ) , .A2( u2_u0_u6_n93 ) );
  NAND4_X1 u2_u0_u6_U79 (.ZN( u2_out0_12 ) , .A4( u2_u0_u6_n114 ) , .A3( u2_u0_u6_n115 ) , .A2( u2_u0_u6_n116 ) , .A1( u2_u0_u6_n117 ) );
  OAI21_X1 u2_u0_u6_U8 (.A( u2_u0_u6_n159 ) , .B1( u2_u0_u6_n169 ) , .B2( u2_u0_u6_n173 ) , .ZN( u2_u0_u6_n90 ) );
  OAI22_X1 u2_u0_u6_U80 (.B2( u2_u0_u6_n111 ) , .ZN( u2_u0_u6_n116 ) , .B1( u2_u0_u6_n126 ) , .A2( u2_u0_u6_n164 ) , .A1( u2_u0_u6_n167 ) );
  OAI21_X1 u2_u0_u6_U81 (.A( u2_u0_u6_n108 ) , .ZN( u2_u0_u6_n117 ) , .B2( u2_u0_u6_n141 ) , .B1( u2_u0_u6_n163 ) );
  OAI211_X1 u2_u0_u6_U82 (.ZN( u2_out0_7 ) , .B( u2_u0_u6_n153 ) , .C2( u2_u0_u6_n154 ) , .C1( u2_u0_u6_n155 ) , .A( u2_u0_u6_n174 ) );
  NOR3_X1 u2_u0_u6_U83 (.A1( u2_u0_u6_n141 ) , .ZN( u2_u0_u6_n154 ) , .A3( u2_u0_u6_n164 ) , .A2( u2_u0_u6_n171 ) );
  AOI211_X1 u2_u0_u6_U84 (.B( u2_u0_u6_n149 ) , .A( u2_u0_u6_n150 ) , .C2( u2_u0_u6_n151 ) , .C1( u2_u0_u6_n152 ) , .ZN( u2_u0_u6_n153 ) );
  OAI211_X1 u2_u0_u6_U85 (.ZN( u2_out0_22 ) , .B( u2_u0_u6_n137 ) , .A( u2_u0_u6_n138 ) , .C2( u2_u0_u6_n139 ) , .C1( u2_u0_u6_n140 ) );
  AOI22_X1 u2_u0_u6_U86 (.B1( u2_u0_u6_n124 ) , .A2( u2_u0_u6_n125 ) , .A1( u2_u0_u6_n126 ) , .ZN( u2_u0_u6_n138 ) , .B2( u2_u0_u6_n161 ) );
  AND4_X1 u2_u0_u6_U87 (.A3( u2_u0_u6_n119 ) , .A1( u2_u0_u6_n120 ) , .A4( u2_u0_u6_n129 ) , .ZN( u2_u0_u6_n140 ) , .A2( u2_u0_u6_n143 ) );
  NAND3_X1 u2_u0_u6_U88 (.A2( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n125 ) , .A1( u2_u0_u6_n130 ) , .A3( u2_u0_u6_n131 ) );
  NAND3_X1 u2_u0_u6_U89 (.A3( u2_u0_u6_n133 ) , .ZN( u2_u0_u6_n141 ) , .A1( u2_u0_u6_n145 ) , .A2( u2_u0_u6_n148 ) );
  INV_X1 u2_u0_u6_U9 (.ZN( u2_u0_u6_n172 ) , .A( u2_u0_u6_n88 ) );
  NAND3_X1 u2_u0_u6_U90 (.ZN( u2_u0_u6_n101 ) , .A3( u2_u0_u6_n107 ) , .A2( u2_u0_u6_n121 ) , .A1( u2_u0_u6_n127 ) );
  NAND3_X1 u2_u0_u6_U91 (.ZN( u2_u0_u6_n102 ) , .A3( u2_u0_u6_n130 ) , .A2( u2_u0_u6_n145 ) , .A1( u2_u0_u6_n166 ) );
  NAND3_X1 u2_u0_u6_U92 (.A3( u2_u0_u6_n113 ) , .A1( u2_u0_u6_n119 ) , .A2( u2_u0_u6_n123 ) , .ZN( u2_u0_u6_n93 ) );
  NAND3_X1 u2_u0_u6_U93 (.ZN( u2_u0_u6_n142 ) , .A2( u2_u0_u6_n172 ) , .A3( u2_u0_u6_n89 ) , .A1( u2_u0_u6_n90 ) );
  INV_X1 u2_u0_u7_U10 (.A( u2_u0_u7_n133 ) , .ZN( u2_u0_u7_n176 ) );
  OAI221_X1 u2_u0_u7_U11 (.C1( u2_u0_u7_n101 ) , .C2( u2_u0_u7_n147 ) , .ZN( u2_u0_u7_n155 ) , .B2( u2_u0_u7_n162 ) , .A( u2_u0_u7_n91 ) , .B1( u2_u0_u7_n92 ) );
  AND3_X1 u2_u0_u7_U12 (.A3( u2_u0_u7_n110 ) , .A2( u2_u0_u7_n127 ) , .A1( u2_u0_u7_n132 ) , .ZN( u2_u0_u7_n92 ) );
  OAI21_X1 u2_u0_u7_U13 (.A( u2_u0_u7_n161 ) , .B1( u2_u0_u7_n168 ) , .B2( u2_u0_u7_n173 ) , .ZN( u2_u0_u7_n91 ) );
  AOI211_X1 u2_u0_u7_U14 (.A( u2_u0_u7_n117 ) , .ZN( u2_u0_u7_n118 ) , .C2( u2_u0_u7_n126 ) , .C1( u2_u0_u7_n177 ) , .B( u2_u0_u7_n180 ) );
  OAI22_X1 u2_u0_u7_U15 (.B1( u2_u0_u7_n115 ) , .ZN( u2_u0_u7_n117 ) , .A2( u2_u0_u7_n133 ) , .A1( u2_u0_u7_n137 ) , .B2( u2_u0_u7_n162 ) );
  INV_X1 u2_u0_u7_U16 (.A( u2_u0_u7_n116 ) , .ZN( u2_u0_u7_n180 ) );
  NOR3_X1 u2_u0_u7_U17 (.ZN( u2_u0_u7_n115 ) , .A3( u2_u0_u7_n145 ) , .A2( u2_u0_u7_n168 ) , .A1( u2_u0_u7_n169 ) );
  NOR3_X1 u2_u0_u7_U18 (.A2( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n135 ) , .ZN( u2_u0_u7_n136 ) , .A3( u2_u0_u7_n171 ) );
  NOR2_X1 u2_u0_u7_U19 (.A1( u2_u0_u7_n130 ) , .A2( u2_u0_u7_n134 ) , .ZN( u2_u0_u7_n153 ) );
  INV_X1 u2_u0_u7_U20 (.A( u2_u0_u7_n101 ) , .ZN( u2_u0_u7_n165 ) );
  NOR2_X1 u2_u0_u7_U21 (.ZN( u2_u0_u7_n111 ) , .A2( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n169 ) );
  AOI21_X1 u2_u0_u7_U22 (.ZN( u2_u0_u7_n104 ) , .B2( u2_u0_u7_n112 ) , .B1( u2_u0_u7_n127 ) , .A( u2_u0_u7_n164 ) );
  AOI21_X1 u2_u0_u7_U23 (.ZN( u2_u0_u7_n106 ) , .B1( u2_u0_u7_n133 ) , .B2( u2_u0_u7_n146 ) , .A( u2_u0_u7_n162 ) );
  AOI21_X1 u2_u0_u7_U24 (.A( u2_u0_u7_n101 ) , .ZN( u2_u0_u7_n107 ) , .B2( u2_u0_u7_n128 ) , .B1( u2_u0_u7_n175 ) );
  INV_X1 u2_u0_u7_U25 (.A( u2_u0_u7_n138 ) , .ZN( u2_u0_u7_n171 ) );
  INV_X1 u2_u0_u7_U26 (.A( u2_u0_u7_n131 ) , .ZN( u2_u0_u7_n177 ) );
  INV_X1 u2_u0_u7_U27 (.A( u2_u0_u7_n110 ) , .ZN( u2_u0_u7_n174 ) );
  NAND2_X1 u2_u0_u7_U28 (.A1( u2_u0_u7_n129 ) , .A2( u2_u0_u7_n132 ) , .ZN( u2_u0_u7_n149 ) );
  NAND2_X1 u2_u0_u7_U29 (.A1( u2_u0_u7_n113 ) , .A2( u2_u0_u7_n124 ) , .ZN( u2_u0_u7_n130 ) );
  OAI21_X1 u2_u0_u7_U3 (.ZN( u2_u0_u7_n159 ) , .A( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n171 ) , .B1( u2_u0_u7_n174 ) );
  INV_X1 u2_u0_u7_U30 (.A( u2_u0_u7_n112 ) , .ZN( u2_u0_u7_n173 ) );
  INV_X1 u2_u0_u7_U31 (.A( u2_u0_u7_n128 ) , .ZN( u2_u0_u7_n168 ) );
  INV_X1 u2_u0_u7_U32 (.A( u2_u0_u7_n148 ) , .ZN( u2_u0_u7_n169 ) );
  INV_X1 u2_u0_u7_U33 (.A( u2_u0_u7_n127 ) , .ZN( u2_u0_u7_n179 ) );
  NOR2_X1 u2_u0_u7_U34 (.ZN( u2_u0_u7_n101 ) , .A2( u2_u0_u7_n150 ) , .A1( u2_u0_u7_n156 ) );
  AOI211_X1 u2_u0_u7_U35 (.B( u2_u0_u7_n139 ) , .A( u2_u0_u7_n140 ) , .C2( u2_u0_u7_n141 ) , .ZN( u2_u0_u7_n142 ) , .C1( u2_u0_u7_n156 ) );
  NAND4_X1 u2_u0_u7_U36 (.A3( u2_u0_u7_n127 ) , .A2( u2_u0_u7_n128 ) , .A1( u2_u0_u7_n129 ) , .ZN( u2_u0_u7_n141 ) , .A4( u2_u0_u7_n147 ) );
  AOI21_X1 u2_u0_u7_U37 (.A( u2_u0_u7_n137 ) , .B1( u2_u0_u7_n138 ) , .ZN( u2_u0_u7_n139 ) , .B2( u2_u0_u7_n146 ) );
  OAI22_X1 u2_u0_u7_U38 (.B1( u2_u0_u7_n136 ) , .ZN( u2_u0_u7_n140 ) , .A1( u2_u0_u7_n153 ) , .B2( u2_u0_u7_n162 ) , .A2( u2_u0_u7_n164 ) );
  AOI211_X1 u2_u0_u7_U39 (.B( u2_u0_u7_n154 ) , .A( u2_u0_u7_n155 ) , .C1( u2_u0_u7_n156 ) , .ZN( u2_u0_u7_n157 ) , .C2( u2_u0_u7_n172 ) );
  INV_X1 u2_u0_u7_U4 (.A( u2_u0_u7_n111 ) , .ZN( u2_u0_u7_n170 ) );
  INV_X1 u2_u0_u7_U40 (.A( u2_u0_u7_n153 ) , .ZN( u2_u0_u7_n172 ) );
  INV_X1 u2_u0_u7_U41 (.A( u2_u0_u7_n125 ) , .ZN( u2_u0_u7_n161 ) );
  NAND2_X1 u2_u0_u7_U42 (.A2( u2_u0_u7_n102 ) , .A1( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n133 ) );
  NAND2_X1 u2_u0_u7_U43 (.A1( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n127 ) , .A2( u2_u0_u7_n99 ) );
  AOI21_X1 u2_u0_u7_U44 (.ZN( u2_u0_u7_n123 ) , .B1( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n177 ) , .A( u2_u0_u7_n97 ) );
  AOI21_X1 u2_u0_u7_U45 (.B2( u2_u0_u7_n113 ) , .B1( u2_u0_u7_n124 ) , .A( u2_u0_u7_n125 ) , .ZN( u2_u0_u7_n97 ) );
  INV_X1 u2_u0_u7_U46 (.A( u2_u0_u7_n152 ) , .ZN( u2_u0_u7_n162 ) );
  AND2_X1 u2_u0_u7_U47 (.ZN( u2_u0_u7_n145 ) , .A2( u2_u0_u7_n98 ) , .A1( u2_u0_u7_n99 ) );
  NOR2_X1 u2_u0_u7_U48 (.ZN( u2_u0_u7_n137 ) , .A1( u2_u0_u7_n150 ) , .A2( u2_u0_u7_n161 ) );
  AOI21_X1 u2_u0_u7_U49 (.ZN( u2_u0_u7_n105 ) , .B2( u2_u0_u7_n110 ) , .A( u2_u0_u7_n125 ) , .B1( u2_u0_u7_n147 ) );
  INV_X1 u2_u0_u7_U5 (.A( u2_u0_u7_n154 ) , .ZN( u2_u0_u7_n178 ) );
  NAND2_X1 u2_u0_u7_U50 (.A2( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n147 ) , .A1( u2_u0_u7_n93 ) );
  NAND2_X1 u2_u0_u7_U51 (.ZN( u2_u0_u7_n146 ) , .A1( u2_u0_u7_n95 ) , .A2( u2_u0_u7_n98 ) );
  OR2_X1 u2_u0_u7_U52 (.ZN( u2_u0_u7_n126 ) , .A2( u2_u0_u7_n152 ) , .A1( u2_u0_u7_n156 ) );
  NAND2_X1 u2_u0_u7_U53 (.ZN( u2_u0_u7_n112 ) , .A2( u2_u0_u7_n96 ) , .A1( u2_u0_u7_n99 ) );
  NAND2_X1 u2_u0_u7_U54 (.A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n128 ) , .A1( u2_u0_u7_n98 ) );
  NAND2_X1 u2_u0_u7_U55 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n113 ) , .A2( u2_u0_u7_n93 ) );
  NAND2_X1 u2_u0_u7_U56 (.ZN( u2_u0_u7_n110 ) , .A1( u2_u0_u7_n95 ) , .A2( u2_u0_u7_n96 ) );
  INV_X1 u2_u0_u7_U57 (.A( u2_u0_u7_n150 ) , .ZN( u2_u0_u7_n164 ) );
  AND2_X1 u2_u0_u7_U58 (.ZN( u2_u0_u7_n134 ) , .A1( u2_u0_u7_n93 ) , .A2( u2_u0_u7_n98 ) );
  NAND2_X1 u2_u0_u7_U59 (.A2( u2_u0_u7_n103 ) , .ZN( u2_u0_u7_n131 ) , .A1( u2_u0_u7_n95 ) );
  INV_X1 u2_u0_u7_U6 (.A( u2_u0_u7_n149 ) , .ZN( u2_u0_u7_n175 ) );
  NAND2_X1 u2_u0_u7_U60 (.A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n124 ) , .A1( u2_u0_u7_n96 ) );
  NAND2_X1 u2_u0_u7_U61 (.A1( u2_u0_u7_n100 ) , .A2( u2_u0_u7_n102 ) , .ZN( u2_u0_u7_n129 ) );
  NAND2_X1 u2_u0_u7_U62 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n138 ) , .A2( u2_u0_u7_n99 ) );
  NAND2_X1 u2_u0_u7_U63 (.ZN( u2_u0_u7_n132 ) , .A1( u2_u0_u7_n93 ) , .A2( u2_u0_u7_n96 ) );
  NAND2_X1 u2_u0_u7_U64 (.A1( u2_u0_u7_n100 ) , .ZN( u2_u0_u7_n148 ) , .A2( u2_u0_u7_n95 ) );
  AOI22_X1 u2_u0_u7_U65 (.A2( u2_u0_u7_n114 ) , .ZN( u2_u0_u7_n119 ) , .B1( u2_u0_u7_n130 ) , .A1( u2_u0_u7_n156 ) , .B2( u2_u0_u7_n165 ) );
  NAND2_X1 u2_u0_u7_U66 (.A2( u2_u0_u7_n112 ) , .ZN( u2_u0_u7_n114 ) , .A1( u2_u0_u7_n175 ) );
  NOR2_X1 u2_u0_u7_U67 (.A2( u2_u0_X_47 ) , .ZN( u2_u0_u7_n150 ) , .A1( u2_u0_u7_n163 ) );
  NOR2_X1 u2_u0_u7_U68 (.A2( u2_u0_X_48 ) , .A1( u2_u0_u7_n166 ) , .ZN( u2_u0_u7_n95 ) );
  NOR2_X1 u2_u0_u7_U69 (.A2( u2_u0_X_45 ) , .A1( u2_u0_X_48 ) , .ZN( u2_u0_u7_n99 ) );
  AOI211_X1 u2_u0_u7_U7 (.ZN( u2_u0_u7_n116 ) , .A( u2_u0_u7_n155 ) , .C1( u2_u0_u7_n161 ) , .C2( u2_u0_u7_n171 ) , .B( u2_u0_u7_n94 ) );
  NOR2_X1 u2_u0_u7_U70 (.A2( u2_u0_X_44 ) , .A1( u2_u0_u7_n167 ) , .ZN( u2_u0_u7_n98 ) );
  NOR2_X1 u2_u0_u7_U71 (.A2( u2_u0_X_46 ) , .A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n152 ) );
  AND2_X1 u2_u0_u7_U72 (.A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n156 ) , .A2( u2_u0_u7_n163 ) );
  NAND2_X1 u2_u0_u7_U73 (.A2( u2_u0_X_46 ) , .A1( u2_u0_X_47 ) , .ZN( u2_u0_u7_n125 ) );
  AND2_X1 u2_u0_u7_U74 (.A2( u2_u0_X_45 ) , .A1( u2_u0_X_48 ) , .ZN( u2_u0_u7_n102 ) );
  AND2_X1 u2_u0_u7_U75 (.A2( u2_u0_X_43 ) , .A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n96 ) );
  AND2_X1 u2_u0_u7_U76 (.A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n100 ) , .A2( u2_u0_u7_n167 ) );
  AND2_X1 u2_u0_u7_U77 (.A1( u2_u0_X_48 ) , .A2( u2_u0_u7_n166 ) , .ZN( u2_u0_u7_n93 ) );
  INV_X1 u2_u0_u7_U78 (.A( u2_u0_X_46 ) , .ZN( u2_u0_u7_n163 ) );
  INV_X1 u2_u0_u7_U79 (.A( u2_u0_X_45 ) , .ZN( u2_u0_u7_n166 ) );
  OAI222_X1 u2_u0_u7_U8 (.C2( u2_u0_u7_n101 ) , .B2( u2_u0_u7_n111 ) , .A1( u2_u0_u7_n113 ) , .C1( u2_u0_u7_n146 ) , .A2( u2_u0_u7_n162 ) , .B1( u2_u0_u7_n164 ) , .ZN( u2_u0_u7_n94 ) );
  OAI21_X1 u2_u0_u7_U80 (.B1( u2_u0_u7_n145 ) , .ZN( u2_u0_u7_n160 ) , .A( u2_u0_u7_n161 ) , .B2( u2_u0_u7_n177 ) );
  AOI22_X1 u2_u0_u7_U81 (.B2( u2_u0_u7_n149 ) , .B1( u2_u0_u7_n150 ) , .A2( u2_u0_u7_n151 ) , .A1( u2_u0_u7_n152 ) , .ZN( u2_u0_u7_n158 ) );
  NAND4_X1 u2_u0_u7_U82 (.ZN( u2_out0_27 ) , .A4( u2_u0_u7_n118 ) , .A3( u2_u0_u7_n119 ) , .A2( u2_u0_u7_n120 ) , .A1( u2_u0_u7_n121 ) );
  OAI21_X1 u2_u0_u7_U83 (.ZN( u2_u0_u7_n121 ) , .B2( u2_u0_u7_n145 ) , .A( u2_u0_u7_n150 ) , .B1( u2_u0_u7_n174 ) );
  OAI21_X1 u2_u0_u7_U84 (.ZN( u2_u0_u7_n120 ) , .A( u2_u0_u7_n161 ) , .B2( u2_u0_u7_n170 ) , .B1( u2_u0_u7_n179 ) );
  NAND4_X1 u2_u0_u7_U85 (.ZN( u2_out0_15 ) , .A4( u2_u0_u7_n142 ) , .A3( u2_u0_u7_n143 ) , .A2( u2_u0_u7_n144 ) , .A1( u2_u0_u7_n178 ) );
  OR2_X1 u2_u0_u7_U86 (.A2( u2_u0_u7_n125 ) , .A1( u2_u0_u7_n129 ) , .ZN( u2_u0_u7_n144 ) );
  AOI22_X1 u2_u0_u7_U87 (.A2( u2_u0_u7_n126 ) , .ZN( u2_u0_u7_n143 ) , .B2( u2_u0_u7_n165 ) , .B1( u2_u0_u7_n173 ) , .A1( u2_u0_u7_n174 ) );
  NAND4_X1 u2_u0_u7_U88 (.ZN( u2_out0_5 ) , .A4( u2_u0_u7_n108 ) , .A3( u2_u0_u7_n109 ) , .A1( u2_u0_u7_n116 ) , .A2( u2_u0_u7_n123 ) );
  AOI22_X1 u2_u0_u7_U89 (.ZN( u2_u0_u7_n109 ) , .A2( u2_u0_u7_n126 ) , .B2( u2_u0_u7_n145 ) , .B1( u2_u0_u7_n156 ) , .A1( u2_u0_u7_n171 ) );
  AOI222_X1 u2_u0_u7_U9 (.ZN( u2_u0_u7_n122 ) , .C2( u2_u0_u7_n126 ) , .C1( u2_u0_u7_n145 ) , .B1( u2_u0_u7_n161 ) , .A2( u2_u0_u7_n165 ) , .B2( u2_u0_u7_n170 ) , .A1( u2_u0_u7_n176 ) );
  NOR4_X1 u2_u0_u7_U90 (.A4( u2_u0_u7_n104 ) , .A3( u2_u0_u7_n105 ) , .A2( u2_u0_u7_n106 ) , .A1( u2_u0_u7_n107 ) , .ZN( u2_u0_u7_n108 ) );
  NAND4_X1 u2_u0_u7_U91 (.ZN( u2_out0_21 ) , .A4( u2_u0_u7_n157 ) , .A3( u2_u0_u7_n158 ) , .A2( u2_u0_u7_n159 ) , .A1( u2_u0_u7_n160 ) );
  OAI211_X1 u2_u0_u7_U92 (.B( u2_u0_u7_n122 ) , .A( u2_u0_u7_n123 ) , .C2( u2_u0_u7_n124 ) , .ZN( u2_u0_u7_n154 ) , .C1( u2_u0_u7_n162 ) );
  NOR2_X1 u2_u0_u7_U93 (.A2( u2_u0_X_43 ) , .A1( u2_u0_X_44 ) , .ZN( u2_u0_u7_n103 ) );
  INV_X1 u2_u0_u7_U94 (.A( u2_u0_X_43 ) , .ZN( u2_u0_u7_n167 ) );
  NAND3_X1 u2_u0_u7_U95 (.A3( u2_u0_u7_n146 ) , .A2( u2_u0_u7_n147 ) , .A1( u2_u0_u7_n148 ) , .ZN( u2_u0_u7_n151 ) );
  NAND3_X1 u2_u0_u7_U96 (.A3( u2_u0_u7_n131 ) , .A2( u2_u0_u7_n132 ) , .A1( u2_u0_u7_n133 ) , .ZN( u2_u0_u7_n135 ) );
  XOR2_X1 u2_u11_U1 (.B( u2_K12_9 ) , .A( u2_R10_6 ) , .Z( u2_u11_X_9 ) );
  XOR2_X1 u2_u11_U16 (.B( u2_K12_3 ) , .A( u2_R10_2 ) , .Z( u2_u11_X_3 ) );
  XOR2_X1 u2_u11_U2 (.B( u2_K12_8 ) , .A( u2_R10_5 ) , .Z( u2_u11_X_8 ) );
  XOR2_X1 u2_u11_U27 (.B( u2_K12_2 ) , .A( u2_R10_1 ) , .Z( u2_u11_X_2 ) );
  XOR2_X1 u2_u11_U3 (.B( u2_K12_7 ) , .A( u2_R10_4 ) , .Z( u2_u11_X_7 ) );
  XOR2_X1 u2_u11_U38 (.B( u2_K12_1 ) , .A( u2_R10_32 ) , .Z( u2_u11_X_1 ) );
  XOR2_X1 u2_u11_U4 (.B( u2_K12_6 ) , .A( u2_R10_5 ) , .Z( u2_u11_X_6 ) );
  XOR2_X1 u2_u11_U46 (.B( u2_K12_12 ) , .A( u2_R10_9 ) , .Z( u2_u11_X_12 ) );
  XOR2_X1 u2_u11_U47 (.B( u2_K12_11 ) , .A( u2_R10_8 ) , .Z( u2_u11_X_11 ) );
  XOR2_X1 u2_u11_U48 (.B( u2_K12_10 ) , .A( u2_R10_7 ) , .Z( u2_u11_X_10 ) );
  XOR2_X1 u2_u11_U5 (.B( u2_K12_5 ) , .A( u2_R10_4 ) , .Z( u2_u11_X_5 ) );
  XOR2_X1 u2_u11_U6 (.B( u2_K12_4 ) , .A( u2_R10_3 ) , .Z( u2_u11_X_4 ) );
  NAND2_X1 u2_u11_u0_U10 (.ZN( u2_u11_u0_n113 ) , .A1( u2_u11_u0_n139 ) , .A2( u2_u11_u0_n149 ) );
  AND3_X1 u2_u11_u0_U11 (.A2( u2_u11_u0_n112 ) , .ZN( u2_u11_u0_n127 ) , .A3( u2_u11_u0_n130 ) , .A1( u2_u11_u0_n148 ) );
  AND2_X1 u2_u11_u0_U12 (.ZN( u2_u11_u0_n107 ) , .A1( u2_u11_u0_n130 ) , .A2( u2_u11_u0_n140 ) );
  AND2_X1 u2_u11_u0_U13 (.A2( u2_u11_u0_n129 ) , .A1( u2_u11_u0_n130 ) , .ZN( u2_u11_u0_n151 ) );
  AND2_X1 u2_u11_u0_U14 (.A1( u2_u11_u0_n108 ) , .A2( u2_u11_u0_n125 ) , .ZN( u2_u11_u0_n145 ) );
  INV_X1 u2_u11_u0_U15 (.A( u2_u11_u0_n143 ) , .ZN( u2_u11_u0_n173 ) );
  NOR2_X1 u2_u11_u0_U16 (.A2( u2_u11_u0_n136 ) , .ZN( u2_u11_u0_n147 ) , .A1( u2_u11_u0_n160 ) );
  OAI22_X1 u2_u11_u0_U17 (.B1( u2_u11_u0_n125 ) , .ZN( u2_u11_u0_n126 ) , .A1( u2_u11_u0_n138 ) , .A2( u2_u11_u0_n146 ) , .B2( u2_u11_u0_n147 ) );
  OAI22_X1 u2_u11_u0_U18 (.B1( u2_u11_u0_n131 ) , .A1( u2_u11_u0_n144 ) , .B2( u2_u11_u0_n147 ) , .A2( u2_u11_u0_n90 ) , .ZN( u2_u11_u0_n91 ) );
  AND3_X1 u2_u11_u0_U19 (.A3( u2_u11_u0_n121 ) , .A2( u2_u11_u0_n125 ) , .A1( u2_u11_u0_n148 ) , .ZN( u2_u11_u0_n90 ) );
  NOR2_X1 u2_u11_u0_U20 (.A1( u2_u11_u0_n163 ) , .A2( u2_u11_u0_n164 ) , .ZN( u2_u11_u0_n95 ) );
  NAND2_X1 u2_u11_u0_U21 (.A1( u2_u11_u0_n101 ) , .A2( u2_u11_u0_n102 ) , .ZN( u2_u11_u0_n150 ) );
  AOI22_X1 u2_u11_u0_U22 (.B2( u2_u11_u0_n109 ) , .A2( u2_u11_u0_n110 ) , .ZN( u2_u11_u0_n111 ) , .B1( u2_u11_u0_n118 ) , .A1( u2_u11_u0_n160 ) );
  NAND2_X1 u2_u11_u0_U23 (.A1( u2_u11_u0_n100 ) , .A2( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n125 ) );
  INV_X1 u2_u11_u0_U24 (.A( u2_u11_u0_n136 ) , .ZN( u2_u11_u0_n161 ) );
  INV_X1 u2_u11_u0_U25 (.A( u2_u11_u0_n118 ) , .ZN( u2_u11_u0_n158 ) );
  NAND2_X1 u2_u11_u0_U26 (.A2( u2_u11_u0_n100 ) , .A1( u2_u11_u0_n101 ) , .ZN( u2_u11_u0_n139 ) );
  NAND2_X1 u2_u11_u0_U27 (.A2( u2_u11_u0_n100 ) , .ZN( u2_u11_u0_n131 ) , .A1( u2_u11_u0_n92 ) );
  NAND2_X1 u2_u11_u0_U28 (.ZN( u2_u11_u0_n108 ) , .A1( u2_u11_u0_n92 ) , .A2( u2_u11_u0_n94 ) );
  AOI21_X1 u2_u11_u0_U29 (.B1( u2_u11_u0_n127 ) , .B2( u2_u11_u0_n129 ) , .A( u2_u11_u0_n138 ) , .ZN( u2_u11_u0_n96 ) );
  INV_X1 u2_u11_u0_U3 (.A( u2_u11_u0_n113 ) , .ZN( u2_u11_u0_n166 ) );
  AOI21_X1 u2_u11_u0_U30 (.ZN( u2_u11_u0_n104 ) , .B1( u2_u11_u0_n107 ) , .B2( u2_u11_u0_n141 ) , .A( u2_u11_u0_n144 ) );
  NAND2_X1 u2_u11_u0_U31 (.A2( u2_u11_u0_n102 ) , .ZN( u2_u11_u0_n114 ) , .A1( u2_u11_u0_n92 ) );
  NAND2_X1 u2_u11_u0_U32 (.A1( u2_u11_u0_n101 ) , .ZN( u2_u11_u0_n130 ) , .A2( u2_u11_u0_n94 ) );
  NOR2_X1 u2_u11_u0_U33 (.A1( u2_u11_u0_n120 ) , .ZN( u2_u11_u0_n143 ) , .A2( u2_u11_u0_n167 ) );
  OAI221_X1 u2_u11_u0_U34 (.C1( u2_u11_u0_n112 ) , .ZN( u2_u11_u0_n120 ) , .B1( u2_u11_u0_n138 ) , .B2( u2_u11_u0_n141 ) , .C2( u2_u11_u0_n147 ) , .A( u2_u11_u0_n172 ) );
  AOI211_X1 u2_u11_u0_U35 (.B( u2_u11_u0_n115 ) , .A( u2_u11_u0_n116 ) , .C2( u2_u11_u0_n117 ) , .C1( u2_u11_u0_n118 ) , .ZN( u2_u11_u0_n119 ) );
  NAND2_X1 u2_u11_u0_U36 (.A2( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n140 ) , .A1( u2_u11_u0_n94 ) );
  INV_X1 u2_u11_u0_U37 (.A( u2_u11_u0_n138 ) , .ZN( u2_u11_u0_n160 ) );
  NAND2_X1 u2_u11_u0_U38 (.A2( u2_u11_u0_n102 ) , .A1( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n149 ) );
  NAND2_X1 u2_u11_u0_U39 (.A2( u2_u11_u0_n101 ) , .ZN( u2_u11_u0_n121 ) , .A1( u2_u11_u0_n93 ) );
  AOI21_X1 u2_u11_u0_U4 (.B1( u2_u11_u0_n114 ) , .ZN( u2_u11_u0_n115 ) , .B2( u2_u11_u0_n129 ) , .A( u2_u11_u0_n161 ) );
  NAND2_X1 u2_u11_u0_U40 (.ZN( u2_u11_u0_n112 ) , .A2( u2_u11_u0_n92 ) , .A1( u2_u11_u0_n93 ) );
  INV_X1 u2_u11_u0_U41 (.ZN( u2_u11_u0_n172 ) , .A( u2_u11_u0_n88 ) );
  OAI222_X1 u2_u11_u0_U42 (.C1( u2_u11_u0_n108 ) , .A1( u2_u11_u0_n125 ) , .B2( u2_u11_u0_n128 ) , .B1( u2_u11_u0_n144 ) , .A2( u2_u11_u0_n158 ) , .C2( u2_u11_u0_n161 ) , .ZN( u2_u11_u0_n88 ) );
  AOI21_X1 u2_u11_u0_U43 (.B1( u2_u11_u0_n103 ) , .ZN( u2_u11_u0_n132 ) , .A( u2_u11_u0_n165 ) , .B2( u2_u11_u0_n93 ) );
  OR3_X1 u2_u11_u0_U44 (.A3( u2_u11_u0_n152 ) , .A2( u2_u11_u0_n153 ) , .A1( u2_u11_u0_n154 ) , .ZN( u2_u11_u0_n155 ) );
  AOI21_X1 u2_u11_u0_U45 (.A( u2_u11_u0_n144 ) , .B2( u2_u11_u0_n145 ) , .B1( u2_u11_u0_n146 ) , .ZN( u2_u11_u0_n154 ) );
  AOI21_X1 u2_u11_u0_U46 (.B2( u2_u11_u0_n150 ) , .B1( u2_u11_u0_n151 ) , .ZN( u2_u11_u0_n152 ) , .A( u2_u11_u0_n158 ) );
  AOI21_X1 u2_u11_u0_U47 (.A( u2_u11_u0_n147 ) , .B2( u2_u11_u0_n148 ) , .B1( u2_u11_u0_n149 ) , .ZN( u2_u11_u0_n153 ) );
  INV_X1 u2_u11_u0_U48 (.ZN( u2_u11_u0_n171 ) , .A( u2_u11_u0_n99 ) );
  OAI211_X1 u2_u11_u0_U49 (.C2( u2_u11_u0_n140 ) , .C1( u2_u11_u0_n161 ) , .A( u2_u11_u0_n169 ) , .B( u2_u11_u0_n98 ) , .ZN( u2_u11_u0_n99 ) );
  AOI21_X1 u2_u11_u0_U5 (.B2( u2_u11_u0_n131 ) , .ZN( u2_u11_u0_n134 ) , .B1( u2_u11_u0_n151 ) , .A( u2_u11_u0_n158 ) );
  AOI211_X1 u2_u11_u0_U50 (.C1( u2_u11_u0_n118 ) , .A( u2_u11_u0_n123 ) , .B( u2_u11_u0_n96 ) , .C2( u2_u11_u0_n97 ) , .ZN( u2_u11_u0_n98 ) );
  INV_X1 u2_u11_u0_U51 (.ZN( u2_u11_u0_n169 ) , .A( u2_u11_u0_n91 ) );
  NOR2_X1 u2_u11_u0_U52 (.A2( u2_u11_X_2 ) , .ZN( u2_u11_u0_n103 ) , .A1( u2_u11_u0_n164 ) );
  NOR2_X1 u2_u11_u0_U53 (.A2( u2_u11_X_4 ) , .A1( u2_u11_X_5 ) , .ZN( u2_u11_u0_n118 ) );
  NOR2_X1 u2_u11_u0_U54 (.A2( u2_u11_X_3 ) , .A1( u2_u11_X_6 ) , .ZN( u2_u11_u0_n94 ) );
  NAND2_X1 u2_u11_u0_U55 (.A2( u2_u11_X_4 ) , .A1( u2_u11_X_5 ) , .ZN( u2_u11_u0_n144 ) );
  NOR2_X1 u2_u11_u0_U56 (.A2( u2_u11_X_5 ) , .ZN( u2_u11_u0_n136 ) , .A1( u2_u11_u0_n159 ) );
  NAND2_X1 u2_u11_u0_U57 (.A1( u2_u11_X_5 ) , .ZN( u2_u11_u0_n138 ) , .A2( u2_u11_u0_n159 ) );
  AND2_X1 u2_u11_u0_U58 (.A2( u2_u11_X_3 ) , .A1( u2_u11_X_6 ) , .ZN( u2_u11_u0_n102 ) );
  AND2_X1 u2_u11_u0_U59 (.A1( u2_u11_X_6 ) , .A2( u2_u11_u0_n162 ) , .ZN( u2_u11_u0_n93 ) );
  NOR2_X1 u2_u11_u0_U6 (.A1( u2_u11_u0_n108 ) , .ZN( u2_u11_u0_n123 ) , .A2( u2_u11_u0_n158 ) );
  INV_X1 u2_u11_u0_U60 (.A( u2_u11_X_4 ) , .ZN( u2_u11_u0_n159 ) );
  INV_X1 u2_u11_u0_U61 (.A( u2_u11_X_2 ) , .ZN( u2_u11_u0_n163 ) );
  INV_X1 u2_u11_u0_U62 (.A( u2_u11_u0_n126 ) , .ZN( u2_u11_u0_n168 ) );
  AOI211_X1 u2_u11_u0_U63 (.B( u2_u11_u0_n133 ) , .A( u2_u11_u0_n134 ) , .C2( u2_u11_u0_n135 ) , .C1( u2_u11_u0_n136 ) , .ZN( u2_u11_u0_n137 ) );
  OR4_X1 u2_u11_u0_U64 (.ZN( u2_out11_17 ) , .A4( u2_u11_u0_n122 ) , .A2( u2_u11_u0_n123 ) , .A1( u2_u11_u0_n124 ) , .A3( u2_u11_u0_n170 ) );
  AOI21_X1 u2_u11_u0_U65 (.B2( u2_u11_u0_n107 ) , .ZN( u2_u11_u0_n124 ) , .B1( u2_u11_u0_n128 ) , .A( u2_u11_u0_n161 ) );
  INV_X1 u2_u11_u0_U66 (.A( u2_u11_u0_n111 ) , .ZN( u2_u11_u0_n170 ) );
  OR4_X1 u2_u11_u0_U67 (.ZN( u2_out11_31 ) , .A4( u2_u11_u0_n155 ) , .A2( u2_u11_u0_n156 ) , .A1( u2_u11_u0_n157 ) , .A3( u2_u11_u0_n173 ) );
  AOI21_X1 u2_u11_u0_U68 (.A( u2_u11_u0_n138 ) , .B2( u2_u11_u0_n139 ) , .B1( u2_u11_u0_n140 ) , .ZN( u2_u11_u0_n157 ) );
  INV_X1 u2_u11_u0_U69 (.ZN( u2_u11_u0_n174 ) , .A( u2_u11_u0_n89 ) );
  OAI21_X1 u2_u11_u0_U7 (.B1( u2_u11_u0_n150 ) , .B2( u2_u11_u0_n158 ) , .A( u2_u11_u0_n172 ) , .ZN( u2_u11_u0_n89 ) );
  AOI211_X1 u2_u11_u0_U70 (.B( u2_u11_u0_n104 ) , .A( u2_u11_u0_n105 ) , .ZN( u2_u11_u0_n106 ) , .C2( u2_u11_u0_n113 ) , .C1( u2_u11_u0_n160 ) );
  INV_X1 u2_u11_u0_U71 (.A( u2_u11_u0_n142 ) , .ZN( u2_u11_u0_n165 ) );
  AOI21_X1 u2_u11_u0_U72 (.ZN( u2_u11_u0_n116 ) , .B2( u2_u11_u0_n142 ) , .A( u2_u11_u0_n144 ) , .B1( u2_u11_u0_n166 ) );
  AOI21_X1 u2_u11_u0_U73 (.B2( u2_u11_u0_n141 ) , .B1( u2_u11_u0_n142 ) , .ZN( u2_u11_u0_n156 ) , .A( u2_u11_u0_n161 ) );
  OAI221_X1 u2_u11_u0_U74 (.C1( u2_u11_u0_n121 ) , .ZN( u2_u11_u0_n122 ) , .B2( u2_u11_u0_n127 ) , .A( u2_u11_u0_n143 ) , .B1( u2_u11_u0_n144 ) , .C2( u2_u11_u0_n147 ) );
  NOR2_X1 u2_u11_u0_U75 (.A2( u2_u11_X_6 ) , .ZN( u2_u11_u0_n100 ) , .A1( u2_u11_u0_n162 ) );
  INV_X1 u2_u11_u0_U76 (.A( u2_u11_X_3 ) , .ZN( u2_u11_u0_n162 ) );
  AOI21_X1 u2_u11_u0_U77 (.B1( u2_u11_u0_n132 ) , .ZN( u2_u11_u0_n133 ) , .A( u2_u11_u0_n144 ) , .B2( u2_u11_u0_n166 ) );
  OAI22_X1 u2_u11_u0_U78 (.ZN( u2_u11_u0_n105 ) , .A2( u2_u11_u0_n132 ) , .B1( u2_u11_u0_n146 ) , .A1( u2_u11_u0_n147 ) , .B2( u2_u11_u0_n161 ) );
  NAND2_X1 u2_u11_u0_U79 (.ZN( u2_u11_u0_n110 ) , .A2( u2_u11_u0_n132 ) , .A1( u2_u11_u0_n145 ) );
  AND2_X1 u2_u11_u0_U8 (.A1( u2_u11_u0_n114 ) , .A2( u2_u11_u0_n121 ) , .ZN( u2_u11_u0_n146 ) );
  INV_X1 u2_u11_u0_U80 (.A( u2_u11_u0_n119 ) , .ZN( u2_u11_u0_n167 ) );
  NAND2_X1 u2_u11_u0_U81 (.ZN( u2_u11_u0_n148 ) , .A1( u2_u11_u0_n93 ) , .A2( u2_u11_u0_n95 ) );
  NAND2_X1 u2_u11_u0_U82 (.A1( u2_u11_u0_n100 ) , .ZN( u2_u11_u0_n129 ) , .A2( u2_u11_u0_n95 ) );
  NAND2_X1 u2_u11_u0_U83 (.A1( u2_u11_u0_n102 ) , .ZN( u2_u11_u0_n128 ) , .A2( u2_u11_u0_n95 ) );
  NOR2_X1 u2_u11_u0_U84 (.A2( u2_u11_X_1 ) , .A1( u2_u11_X_2 ) , .ZN( u2_u11_u0_n92 ) );
  NAND2_X1 u2_u11_u0_U85 (.ZN( u2_u11_u0_n142 ) , .A1( u2_u11_u0_n94 ) , .A2( u2_u11_u0_n95 ) );
  NOR2_X1 u2_u11_u0_U86 (.A2( u2_u11_X_1 ) , .ZN( u2_u11_u0_n101 ) , .A1( u2_u11_u0_n163 ) );
  INV_X1 u2_u11_u0_U87 (.A( u2_u11_X_1 ) , .ZN( u2_u11_u0_n164 ) );
  NAND3_X1 u2_u11_u0_U88 (.ZN( u2_out11_23 ) , .A3( u2_u11_u0_n137 ) , .A1( u2_u11_u0_n168 ) , .A2( u2_u11_u0_n171 ) );
  NAND3_X1 u2_u11_u0_U89 (.A3( u2_u11_u0_n127 ) , .A2( u2_u11_u0_n128 ) , .ZN( u2_u11_u0_n135 ) , .A1( u2_u11_u0_n150 ) );
  AND2_X1 u2_u11_u0_U9 (.A1( u2_u11_u0_n131 ) , .ZN( u2_u11_u0_n141 ) , .A2( u2_u11_u0_n150 ) );
  NAND3_X1 u2_u11_u0_U90 (.ZN( u2_u11_u0_n117 ) , .A3( u2_u11_u0_n132 ) , .A2( u2_u11_u0_n139 ) , .A1( u2_u11_u0_n148 ) );
  NAND3_X1 u2_u11_u0_U91 (.ZN( u2_u11_u0_n109 ) , .A2( u2_u11_u0_n114 ) , .A3( u2_u11_u0_n140 ) , .A1( u2_u11_u0_n149 ) );
  NAND3_X1 u2_u11_u0_U92 (.ZN( u2_out11_9 ) , .A3( u2_u11_u0_n106 ) , .A2( u2_u11_u0_n171 ) , .A1( u2_u11_u0_n174 ) );
  NAND3_X1 u2_u11_u0_U93 (.A2( u2_u11_u0_n128 ) , .A1( u2_u11_u0_n132 ) , .A3( u2_u11_u0_n146 ) , .ZN( u2_u11_u0_n97 ) );
  NOR2_X1 u2_u11_u1_U10 (.A1( u2_u11_u1_n112 ) , .A2( u2_u11_u1_n116 ) , .ZN( u2_u11_u1_n118 ) );
  NAND3_X1 u2_u11_u1_U100 (.ZN( u2_u11_u1_n113 ) , .A1( u2_u11_u1_n120 ) , .A3( u2_u11_u1_n133 ) , .A2( u2_u11_u1_n155 ) );
  OAI21_X1 u2_u11_u1_U11 (.ZN( u2_u11_u1_n101 ) , .B1( u2_u11_u1_n141 ) , .A( u2_u11_u1_n146 ) , .B2( u2_u11_u1_n183 ) );
  AOI21_X1 u2_u11_u1_U12 (.B2( u2_u11_u1_n155 ) , .B1( u2_u11_u1_n156 ) , .ZN( u2_u11_u1_n157 ) , .A( u2_u11_u1_n174 ) );
  NAND2_X1 u2_u11_u1_U13 (.ZN( u2_u11_u1_n140 ) , .A2( u2_u11_u1_n150 ) , .A1( u2_u11_u1_n155 ) );
  NAND2_X1 u2_u11_u1_U14 (.A1( u2_u11_u1_n131 ) , .ZN( u2_u11_u1_n147 ) , .A2( u2_u11_u1_n153 ) );
  INV_X1 u2_u11_u1_U15 (.A( u2_u11_u1_n139 ) , .ZN( u2_u11_u1_n174 ) );
  OR4_X1 u2_u11_u1_U16 (.A4( u2_u11_u1_n106 ) , .A3( u2_u11_u1_n107 ) , .ZN( u2_u11_u1_n108 ) , .A1( u2_u11_u1_n117 ) , .A2( u2_u11_u1_n184 ) );
  AOI21_X1 u2_u11_u1_U17 (.ZN( u2_u11_u1_n106 ) , .A( u2_u11_u1_n112 ) , .B1( u2_u11_u1_n154 ) , .B2( u2_u11_u1_n156 ) );
  AOI21_X1 u2_u11_u1_U18 (.ZN( u2_u11_u1_n107 ) , .B1( u2_u11_u1_n134 ) , .B2( u2_u11_u1_n149 ) , .A( u2_u11_u1_n174 ) );
  INV_X1 u2_u11_u1_U19 (.A( u2_u11_u1_n101 ) , .ZN( u2_u11_u1_n184 ) );
  INV_X1 u2_u11_u1_U20 (.A( u2_u11_u1_n112 ) , .ZN( u2_u11_u1_n171 ) );
  NAND2_X1 u2_u11_u1_U21 (.ZN( u2_u11_u1_n141 ) , .A1( u2_u11_u1_n153 ) , .A2( u2_u11_u1_n156 ) );
  AND2_X1 u2_u11_u1_U22 (.A1( u2_u11_u1_n123 ) , .ZN( u2_u11_u1_n134 ) , .A2( u2_u11_u1_n161 ) );
  NAND2_X1 u2_u11_u1_U23 (.A2( u2_u11_u1_n115 ) , .A1( u2_u11_u1_n116 ) , .ZN( u2_u11_u1_n148 ) );
  NAND2_X1 u2_u11_u1_U24 (.A2( u2_u11_u1_n133 ) , .A1( u2_u11_u1_n135 ) , .ZN( u2_u11_u1_n159 ) );
  NAND2_X1 u2_u11_u1_U25 (.A2( u2_u11_u1_n115 ) , .A1( u2_u11_u1_n120 ) , .ZN( u2_u11_u1_n132 ) );
  INV_X1 u2_u11_u1_U26 (.A( u2_u11_u1_n154 ) , .ZN( u2_u11_u1_n178 ) );
  INV_X1 u2_u11_u1_U27 (.A( u2_u11_u1_n151 ) , .ZN( u2_u11_u1_n183 ) );
  AND2_X1 u2_u11_u1_U28 (.A1( u2_u11_u1_n129 ) , .A2( u2_u11_u1_n133 ) , .ZN( u2_u11_u1_n149 ) );
  INV_X1 u2_u11_u1_U29 (.A( u2_u11_u1_n131 ) , .ZN( u2_u11_u1_n180 ) );
  INV_X1 u2_u11_u1_U3 (.A( u2_u11_u1_n159 ) , .ZN( u2_u11_u1_n182 ) );
  OAI221_X1 u2_u11_u1_U30 (.A( u2_u11_u1_n119 ) , .C2( u2_u11_u1_n129 ) , .ZN( u2_u11_u1_n138 ) , .B2( u2_u11_u1_n152 ) , .C1( u2_u11_u1_n174 ) , .B1( u2_u11_u1_n187 ) );
  INV_X1 u2_u11_u1_U31 (.A( u2_u11_u1_n148 ) , .ZN( u2_u11_u1_n187 ) );
  AOI211_X1 u2_u11_u1_U32 (.B( u2_u11_u1_n117 ) , .A( u2_u11_u1_n118 ) , .ZN( u2_u11_u1_n119 ) , .C2( u2_u11_u1_n146 ) , .C1( u2_u11_u1_n159 ) );
  NOR2_X1 u2_u11_u1_U33 (.A1( u2_u11_u1_n168 ) , .A2( u2_u11_u1_n176 ) , .ZN( u2_u11_u1_n98 ) );
  AOI211_X1 u2_u11_u1_U34 (.B( u2_u11_u1_n162 ) , .A( u2_u11_u1_n163 ) , .C2( u2_u11_u1_n164 ) , .ZN( u2_u11_u1_n165 ) , .C1( u2_u11_u1_n171 ) );
  AOI21_X1 u2_u11_u1_U35 (.A( u2_u11_u1_n160 ) , .B2( u2_u11_u1_n161 ) , .ZN( u2_u11_u1_n162 ) , .B1( u2_u11_u1_n182 ) );
  OR2_X1 u2_u11_u1_U36 (.A2( u2_u11_u1_n157 ) , .A1( u2_u11_u1_n158 ) , .ZN( u2_u11_u1_n163 ) );
  NAND2_X1 u2_u11_u1_U37 (.A1( u2_u11_u1_n128 ) , .ZN( u2_u11_u1_n146 ) , .A2( u2_u11_u1_n160 ) );
  NAND2_X1 u2_u11_u1_U38 (.A2( u2_u11_u1_n112 ) , .ZN( u2_u11_u1_n139 ) , .A1( u2_u11_u1_n152 ) );
  NAND2_X1 u2_u11_u1_U39 (.A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n156 ) , .A2( u2_u11_u1_n99 ) );
  AOI221_X1 u2_u11_u1_U4 (.A( u2_u11_u1_n138 ) , .C2( u2_u11_u1_n139 ) , .C1( u2_u11_u1_n140 ) , .B2( u2_u11_u1_n141 ) , .ZN( u2_u11_u1_n142 ) , .B1( u2_u11_u1_n175 ) );
  AOI221_X1 u2_u11_u1_U40 (.B1( u2_u11_u1_n140 ) , .ZN( u2_u11_u1_n167 ) , .B2( u2_u11_u1_n172 ) , .C2( u2_u11_u1_n175 ) , .C1( u2_u11_u1_n178 ) , .A( u2_u11_u1_n188 ) );
  INV_X1 u2_u11_u1_U41 (.ZN( u2_u11_u1_n188 ) , .A( u2_u11_u1_n97 ) );
  AOI211_X1 u2_u11_u1_U42 (.A( u2_u11_u1_n118 ) , .C1( u2_u11_u1_n132 ) , .C2( u2_u11_u1_n139 ) , .B( u2_u11_u1_n96 ) , .ZN( u2_u11_u1_n97 ) );
  AOI21_X1 u2_u11_u1_U43 (.B2( u2_u11_u1_n121 ) , .B1( u2_u11_u1_n135 ) , .A( u2_u11_u1_n152 ) , .ZN( u2_u11_u1_n96 ) );
  NOR2_X1 u2_u11_u1_U44 (.ZN( u2_u11_u1_n117 ) , .A1( u2_u11_u1_n121 ) , .A2( u2_u11_u1_n160 ) );
  OAI21_X1 u2_u11_u1_U45 (.B2( u2_u11_u1_n123 ) , .ZN( u2_u11_u1_n145 ) , .B1( u2_u11_u1_n160 ) , .A( u2_u11_u1_n185 ) );
  INV_X1 u2_u11_u1_U46 (.A( u2_u11_u1_n122 ) , .ZN( u2_u11_u1_n185 ) );
  AOI21_X1 u2_u11_u1_U47 (.B2( u2_u11_u1_n120 ) , .B1( u2_u11_u1_n121 ) , .ZN( u2_u11_u1_n122 ) , .A( u2_u11_u1_n128 ) );
  AOI21_X1 u2_u11_u1_U48 (.A( u2_u11_u1_n128 ) , .B2( u2_u11_u1_n129 ) , .ZN( u2_u11_u1_n130 ) , .B1( u2_u11_u1_n150 ) );
  NAND2_X1 u2_u11_u1_U49 (.ZN( u2_u11_u1_n112 ) , .A1( u2_u11_u1_n169 ) , .A2( u2_u11_u1_n170 ) );
  AOI211_X1 u2_u11_u1_U5 (.ZN( u2_u11_u1_n124 ) , .A( u2_u11_u1_n138 ) , .C2( u2_u11_u1_n139 ) , .B( u2_u11_u1_n145 ) , .C1( u2_u11_u1_n147 ) );
  NAND2_X1 u2_u11_u1_U50 (.ZN( u2_u11_u1_n129 ) , .A2( u2_u11_u1_n95 ) , .A1( u2_u11_u1_n98 ) );
  NAND2_X1 u2_u11_u1_U51 (.A1( u2_u11_u1_n102 ) , .ZN( u2_u11_u1_n154 ) , .A2( u2_u11_u1_n99 ) );
  NAND2_X1 u2_u11_u1_U52 (.A2( u2_u11_u1_n100 ) , .ZN( u2_u11_u1_n135 ) , .A1( u2_u11_u1_n99 ) );
  AOI21_X1 u2_u11_u1_U53 (.A( u2_u11_u1_n152 ) , .B2( u2_u11_u1_n153 ) , .B1( u2_u11_u1_n154 ) , .ZN( u2_u11_u1_n158 ) );
  INV_X1 u2_u11_u1_U54 (.A( u2_u11_u1_n160 ) , .ZN( u2_u11_u1_n175 ) );
  NAND2_X1 u2_u11_u1_U55 (.A1( u2_u11_u1_n100 ) , .ZN( u2_u11_u1_n116 ) , .A2( u2_u11_u1_n95 ) );
  NAND2_X1 u2_u11_u1_U56 (.A1( u2_u11_u1_n102 ) , .ZN( u2_u11_u1_n131 ) , .A2( u2_u11_u1_n95 ) );
  NAND2_X1 u2_u11_u1_U57 (.A2( u2_u11_u1_n104 ) , .ZN( u2_u11_u1_n121 ) , .A1( u2_u11_u1_n98 ) );
  NAND2_X1 u2_u11_u1_U58 (.A1( u2_u11_u1_n103 ) , .ZN( u2_u11_u1_n153 ) , .A2( u2_u11_u1_n98 ) );
  NAND2_X1 u2_u11_u1_U59 (.A2( u2_u11_u1_n104 ) , .A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n133 ) );
  AOI22_X1 u2_u11_u1_U6 (.B2( u2_u11_u1_n113 ) , .A2( u2_u11_u1_n114 ) , .ZN( u2_u11_u1_n125 ) , .A1( u2_u11_u1_n171 ) , .B1( u2_u11_u1_n173 ) );
  NAND2_X1 u2_u11_u1_U60 (.ZN( u2_u11_u1_n150 ) , .A2( u2_u11_u1_n98 ) , .A1( u2_u11_u1_n99 ) );
  NAND2_X1 u2_u11_u1_U61 (.A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n155 ) , .A2( u2_u11_u1_n95 ) );
  OAI21_X1 u2_u11_u1_U62 (.ZN( u2_u11_u1_n109 ) , .B1( u2_u11_u1_n129 ) , .B2( u2_u11_u1_n160 ) , .A( u2_u11_u1_n167 ) );
  NAND2_X1 u2_u11_u1_U63 (.A2( u2_u11_u1_n100 ) , .A1( u2_u11_u1_n103 ) , .ZN( u2_u11_u1_n120 ) );
  NAND2_X1 u2_u11_u1_U64 (.A1( u2_u11_u1_n102 ) , .A2( u2_u11_u1_n104 ) , .ZN( u2_u11_u1_n115 ) );
  NAND2_X1 u2_u11_u1_U65 (.A2( u2_u11_u1_n100 ) , .A1( u2_u11_u1_n104 ) , .ZN( u2_u11_u1_n151 ) );
  NAND2_X1 u2_u11_u1_U66 (.A2( u2_u11_u1_n103 ) , .A1( u2_u11_u1_n105 ) , .ZN( u2_u11_u1_n161 ) );
  INV_X1 u2_u11_u1_U67 (.A( u2_u11_u1_n152 ) , .ZN( u2_u11_u1_n173 ) );
  INV_X1 u2_u11_u1_U68 (.A( u2_u11_u1_n128 ) , .ZN( u2_u11_u1_n172 ) );
  NAND2_X1 u2_u11_u1_U69 (.A2( u2_u11_u1_n102 ) , .A1( u2_u11_u1_n103 ) , .ZN( u2_u11_u1_n123 ) );
  NAND2_X1 u2_u11_u1_U7 (.ZN( u2_u11_u1_n114 ) , .A1( u2_u11_u1_n134 ) , .A2( u2_u11_u1_n156 ) );
  NOR2_X1 u2_u11_u1_U70 (.A2( u2_u11_X_7 ) , .A1( u2_u11_X_8 ) , .ZN( u2_u11_u1_n95 ) );
  NOR2_X1 u2_u11_u1_U71 (.A1( u2_u11_X_12 ) , .A2( u2_u11_X_9 ) , .ZN( u2_u11_u1_n100 ) );
  NOR2_X1 u2_u11_u1_U72 (.A2( u2_u11_X_8 ) , .A1( u2_u11_u1_n177 ) , .ZN( u2_u11_u1_n99 ) );
  NOR2_X1 u2_u11_u1_U73 (.A2( u2_u11_X_12 ) , .ZN( u2_u11_u1_n102 ) , .A1( u2_u11_u1_n176 ) );
  NOR2_X1 u2_u11_u1_U74 (.A2( u2_u11_X_9 ) , .ZN( u2_u11_u1_n105 ) , .A1( u2_u11_u1_n168 ) );
  NAND2_X1 u2_u11_u1_U75 (.A1( u2_u11_X_10 ) , .ZN( u2_u11_u1_n160 ) , .A2( u2_u11_u1_n169 ) );
  NAND2_X1 u2_u11_u1_U76 (.A2( u2_u11_X_10 ) , .A1( u2_u11_X_11 ) , .ZN( u2_u11_u1_n152 ) );
  NAND2_X1 u2_u11_u1_U77 (.A1( u2_u11_X_11 ) , .ZN( u2_u11_u1_n128 ) , .A2( u2_u11_u1_n170 ) );
  AND2_X1 u2_u11_u1_U78 (.A2( u2_u11_X_7 ) , .A1( u2_u11_X_8 ) , .ZN( u2_u11_u1_n104 ) );
  AND2_X1 u2_u11_u1_U79 (.A1( u2_u11_X_8 ) , .ZN( u2_u11_u1_n103 ) , .A2( u2_u11_u1_n177 ) );
  AOI22_X1 u2_u11_u1_U8 (.B2( u2_u11_u1_n136 ) , .A2( u2_u11_u1_n137 ) , .ZN( u2_u11_u1_n143 ) , .A1( u2_u11_u1_n171 ) , .B1( u2_u11_u1_n173 ) );
  INV_X1 u2_u11_u1_U80 (.A( u2_u11_X_10 ) , .ZN( u2_u11_u1_n170 ) );
  INV_X1 u2_u11_u1_U81 (.A( u2_u11_X_9 ) , .ZN( u2_u11_u1_n176 ) );
  INV_X1 u2_u11_u1_U82 (.A( u2_u11_X_11 ) , .ZN( u2_u11_u1_n169 ) );
  INV_X1 u2_u11_u1_U83 (.A( u2_u11_X_12 ) , .ZN( u2_u11_u1_n168 ) );
  INV_X1 u2_u11_u1_U84 (.A( u2_u11_X_7 ) , .ZN( u2_u11_u1_n177 ) );
  NAND4_X1 u2_u11_u1_U85 (.ZN( u2_out11_28 ) , .A4( u2_u11_u1_n124 ) , .A3( u2_u11_u1_n125 ) , .A2( u2_u11_u1_n126 ) , .A1( u2_u11_u1_n127 ) );
  OAI21_X1 u2_u11_u1_U86 (.ZN( u2_u11_u1_n127 ) , .B2( u2_u11_u1_n139 ) , .B1( u2_u11_u1_n175 ) , .A( u2_u11_u1_n183 ) );
  OAI21_X1 u2_u11_u1_U87 (.ZN( u2_u11_u1_n126 ) , .B2( u2_u11_u1_n140 ) , .A( u2_u11_u1_n146 ) , .B1( u2_u11_u1_n178 ) );
  NAND4_X1 u2_u11_u1_U88 (.ZN( u2_out11_18 ) , .A4( u2_u11_u1_n165 ) , .A3( u2_u11_u1_n166 ) , .A1( u2_u11_u1_n167 ) , .A2( u2_u11_u1_n186 ) );
  AOI22_X1 u2_u11_u1_U89 (.B2( u2_u11_u1_n146 ) , .B1( u2_u11_u1_n147 ) , .A2( u2_u11_u1_n148 ) , .ZN( u2_u11_u1_n166 ) , .A1( u2_u11_u1_n172 ) );
  INV_X1 u2_u11_u1_U9 (.A( u2_u11_u1_n147 ) , .ZN( u2_u11_u1_n181 ) );
  INV_X1 u2_u11_u1_U90 (.A( u2_u11_u1_n145 ) , .ZN( u2_u11_u1_n186 ) );
  NAND4_X1 u2_u11_u1_U91 (.ZN( u2_out11_2 ) , .A4( u2_u11_u1_n142 ) , .A3( u2_u11_u1_n143 ) , .A2( u2_u11_u1_n144 ) , .A1( u2_u11_u1_n179 ) );
  OAI21_X1 u2_u11_u1_U92 (.B2( u2_u11_u1_n132 ) , .ZN( u2_u11_u1_n144 ) , .A( u2_u11_u1_n146 ) , .B1( u2_u11_u1_n180 ) );
  INV_X1 u2_u11_u1_U93 (.A( u2_u11_u1_n130 ) , .ZN( u2_u11_u1_n179 ) );
  OR4_X1 u2_u11_u1_U94 (.ZN( u2_out11_13 ) , .A4( u2_u11_u1_n108 ) , .A3( u2_u11_u1_n109 ) , .A2( u2_u11_u1_n110 ) , .A1( u2_u11_u1_n111 ) );
  AOI21_X1 u2_u11_u1_U95 (.ZN( u2_u11_u1_n111 ) , .A( u2_u11_u1_n128 ) , .B2( u2_u11_u1_n131 ) , .B1( u2_u11_u1_n135 ) );
  AOI21_X1 u2_u11_u1_U96 (.ZN( u2_u11_u1_n110 ) , .A( u2_u11_u1_n116 ) , .B1( u2_u11_u1_n152 ) , .B2( u2_u11_u1_n160 ) );
  NAND3_X1 u2_u11_u1_U97 (.A3( u2_u11_u1_n149 ) , .A2( u2_u11_u1_n150 ) , .A1( u2_u11_u1_n151 ) , .ZN( u2_u11_u1_n164 ) );
  NAND3_X1 u2_u11_u1_U98 (.A3( u2_u11_u1_n134 ) , .A2( u2_u11_u1_n135 ) , .ZN( u2_u11_u1_n136 ) , .A1( u2_u11_u1_n151 ) );
  NAND3_X1 u2_u11_u1_U99 (.A1( u2_u11_u1_n133 ) , .ZN( u2_u11_u1_n137 ) , .A2( u2_u11_u1_n154 ) , .A3( u2_u11_u1_n181 ) );
  XOR2_X1 u2_u13_U10 (.B( u2_K14_45 ) , .A( u2_R12_30 ) , .Z( u2_u13_X_45 ) );
  XOR2_X1 u2_u13_U11 (.B( u2_K14_44 ) , .A( u2_R12_29 ) , .Z( u2_u13_X_44 ) );
  XOR2_X1 u2_u13_U12 (.B( u2_K14_43 ) , .A( u2_R12_28 ) , .Z( u2_u13_X_43 ) );
  XOR2_X1 u2_u13_U7 (.B( u2_K14_48 ) , .A( u2_R12_1 ) , .Z( u2_u13_X_48 ) );
  XOR2_X1 u2_u13_U8 (.B( u2_K14_47 ) , .A( u2_R12_32 ) , .Z( u2_u13_X_47 ) );
  XOR2_X1 u2_u13_U9 (.B( u2_K14_46 ) , .A( u2_R12_31 ) , .Z( u2_u13_X_46 ) );
  AND3_X1 u2_u13_u7_U10 (.A3( u2_u13_u7_n110 ) , .A2( u2_u13_u7_n127 ) , .A1( u2_u13_u7_n132 ) , .ZN( u2_u13_u7_n92 ) );
  OAI21_X1 u2_u13_u7_U11 (.A( u2_u13_u7_n161 ) , .B1( u2_u13_u7_n168 ) , .B2( u2_u13_u7_n173 ) , .ZN( u2_u13_u7_n91 ) );
  AOI211_X1 u2_u13_u7_U12 (.A( u2_u13_u7_n117 ) , .ZN( u2_u13_u7_n118 ) , .C2( u2_u13_u7_n126 ) , .C1( u2_u13_u7_n177 ) , .B( u2_u13_u7_n180 ) );
  OAI22_X1 u2_u13_u7_U13 (.B1( u2_u13_u7_n115 ) , .ZN( u2_u13_u7_n117 ) , .A2( u2_u13_u7_n133 ) , .A1( u2_u13_u7_n137 ) , .B2( u2_u13_u7_n162 ) );
  INV_X1 u2_u13_u7_U14 (.A( u2_u13_u7_n116 ) , .ZN( u2_u13_u7_n180 ) );
  NOR3_X1 u2_u13_u7_U15 (.ZN( u2_u13_u7_n115 ) , .A3( u2_u13_u7_n145 ) , .A2( u2_u13_u7_n168 ) , .A1( u2_u13_u7_n169 ) );
  OAI211_X1 u2_u13_u7_U16 (.B( u2_u13_u7_n122 ) , .A( u2_u13_u7_n123 ) , .C2( u2_u13_u7_n124 ) , .ZN( u2_u13_u7_n154 ) , .C1( u2_u13_u7_n162 ) );
  AOI222_X1 u2_u13_u7_U17 (.ZN( u2_u13_u7_n122 ) , .C2( u2_u13_u7_n126 ) , .C1( u2_u13_u7_n145 ) , .B1( u2_u13_u7_n161 ) , .A2( u2_u13_u7_n165 ) , .B2( u2_u13_u7_n170 ) , .A1( u2_u13_u7_n176 ) );
  INV_X1 u2_u13_u7_U18 (.A( u2_u13_u7_n133 ) , .ZN( u2_u13_u7_n176 ) );
  NOR3_X1 u2_u13_u7_U19 (.A2( u2_u13_u7_n134 ) , .A1( u2_u13_u7_n135 ) , .ZN( u2_u13_u7_n136 ) , .A3( u2_u13_u7_n171 ) );
  NOR2_X1 u2_u13_u7_U20 (.A1( u2_u13_u7_n130 ) , .A2( u2_u13_u7_n134 ) , .ZN( u2_u13_u7_n153 ) );
  INV_X1 u2_u13_u7_U21 (.A( u2_u13_u7_n101 ) , .ZN( u2_u13_u7_n165 ) );
  NOR2_X1 u2_u13_u7_U22 (.ZN( u2_u13_u7_n111 ) , .A2( u2_u13_u7_n134 ) , .A1( u2_u13_u7_n169 ) );
  AOI21_X1 u2_u13_u7_U23 (.ZN( u2_u13_u7_n104 ) , .B2( u2_u13_u7_n112 ) , .B1( u2_u13_u7_n127 ) , .A( u2_u13_u7_n164 ) );
  AOI21_X1 u2_u13_u7_U24 (.ZN( u2_u13_u7_n106 ) , .B1( u2_u13_u7_n133 ) , .B2( u2_u13_u7_n146 ) , .A( u2_u13_u7_n162 ) );
  AOI21_X1 u2_u13_u7_U25 (.A( u2_u13_u7_n101 ) , .ZN( u2_u13_u7_n107 ) , .B2( u2_u13_u7_n128 ) , .B1( u2_u13_u7_n175 ) );
  INV_X1 u2_u13_u7_U26 (.A( u2_u13_u7_n138 ) , .ZN( u2_u13_u7_n171 ) );
  INV_X1 u2_u13_u7_U27 (.A( u2_u13_u7_n131 ) , .ZN( u2_u13_u7_n177 ) );
  INV_X1 u2_u13_u7_U28 (.A( u2_u13_u7_n110 ) , .ZN( u2_u13_u7_n174 ) );
  NAND2_X1 u2_u13_u7_U29 (.A1( u2_u13_u7_n129 ) , .A2( u2_u13_u7_n132 ) , .ZN( u2_u13_u7_n149 ) );
  OAI21_X1 u2_u13_u7_U3 (.ZN( u2_u13_u7_n159 ) , .A( u2_u13_u7_n165 ) , .B2( u2_u13_u7_n171 ) , .B1( u2_u13_u7_n174 ) );
  NAND2_X1 u2_u13_u7_U30 (.A1( u2_u13_u7_n113 ) , .A2( u2_u13_u7_n124 ) , .ZN( u2_u13_u7_n130 ) );
  INV_X1 u2_u13_u7_U31 (.A( u2_u13_u7_n112 ) , .ZN( u2_u13_u7_n173 ) );
  INV_X1 u2_u13_u7_U32 (.A( u2_u13_u7_n128 ) , .ZN( u2_u13_u7_n168 ) );
  INV_X1 u2_u13_u7_U33 (.A( u2_u13_u7_n148 ) , .ZN( u2_u13_u7_n169 ) );
  INV_X1 u2_u13_u7_U34 (.A( u2_u13_u7_n127 ) , .ZN( u2_u13_u7_n179 ) );
  NOR2_X1 u2_u13_u7_U35 (.ZN( u2_u13_u7_n101 ) , .A2( u2_u13_u7_n150 ) , .A1( u2_u13_u7_n156 ) );
  AOI211_X1 u2_u13_u7_U36 (.B( u2_u13_u7_n154 ) , .A( u2_u13_u7_n155 ) , .C1( u2_u13_u7_n156 ) , .ZN( u2_u13_u7_n157 ) , .C2( u2_u13_u7_n172 ) );
  INV_X1 u2_u13_u7_U37 (.A( u2_u13_u7_n153 ) , .ZN( u2_u13_u7_n172 ) );
  AOI211_X1 u2_u13_u7_U38 (.B( u2_u13_u7_n139 ) , .A( u2_u13_u7_n140 ) , .C2( u2_u13_u7_n141 ) , .ZN( u2_u13_u7_n142 ) , .C1( u2_u13_u7_n156 ) );
  NAND4_X1 u2_u13_u7_U39 (.A3( u2_u13_u7_n127 ) , .A2( u2_u13_u7_n128 ) , .A1( u2_u13_u7_n129 ) , .ZN( u2_u13_u7_n141 ) , .A4( u2_u13_u7_n147 ) );
  INV_X1 u2_u13_u7_U4 (.A( u2_u13_u7_n111 ) , .ZN( u2_u13_u7_n170 ) );
  AOI21_X1 u2_u13_u7_U40 (.A( u2_u13_u7_n137 ) , .B1( u2_u13_u7_n138 ) , .ZN( u2_u13_u7_n139 ) , .B2( u2_u13_u7_n146 ) );
  OAI22_X1 u2_u13_u7_U41 (.B1( u2_u13_u7_n136 ) , .ZN( u2_u13_u7_n140 ) , .A1( u2_u13_u7_n153 ) , .B2( u2_u13_u7_n162 ) , .A2( u2_u13_u7_n164 ) );
  AOI21_X1 u2_u13_u7_U42 (.ZN( u2_u13_u7_n123 ) , .B1( u2_u13_u7_n165 ) , .B2( u2_u13_u7_n177 ) , .A( u2_u13_u7_n97 ) );
  AOI21_X1 u2_u13_u7_U43 (.B2( u2_u13_u7_n113 ) , .B1( u2_u13_u7_n124 ) , .A( u2_u13_u7_n125 ) , .ZN( u2_u13_u7_n97 ) );
  INV_X1 u2_u13_u7_U44 (.A( u2_u13_u7_n125 ) , .ZN( u2_u13_u7_n161 ) );
  INV_X1 u2_u13_u7_U45 (.A( u2_u13_u7_n152 ) , .ZN( u2_u13_u7_n162 ) );
  AOI22_X1 u2_u13_u7_U46 (.A2( u2_u13_u7_n114 ) , .ZN( u2_u13_u7_n119 ) , .B1( u2_u13_u7_n130 ) , .A1( u2_u13_u7_n156 ) , .B2( u2_u13_u7_n165 ) );
  NAND2_X1 u2_u13_u7_U47 (.A2( u2_u13_u7_n112 ) , .ZN( u2_u13_u7_n114 ) , .A1( u2_u13_u7_n175 ) );
  AND2_X1 u2_u13_u7_U48 (.ZN( u2_u13_u7_n145 ) , .A2( u2_u13_u7_n98 ) , .A1( u2_u13_u7_n99 ) );
  NOR2_X1 u2_u13_u7_U49 (.ZN( u2_u13_u7_n137 ) , .A1( u2_u13_u7_n150 ) , .A2( u2_u13_u7_n161 ) );
  INV_X1 u2_u13_u7_U5 (.A( u2_u13_u7_n149 ) , .ZN( u2_u13_u7_n175 ) );
  AOI21_X1 u2_u13_u7_U50 (.ZN( u2_u13_u7_n105 ) , .B2( u2_u13_u7_n110 ) , .A( u2_u13_u7_n125 ) , .B1( u2_u13_u7_n147 ) );
  NAND2_X1 u2_u13_u7_U51 (.ZN( u2_u13_u7_n146 ) , .A1( u2_u13_u7_n95 ) , .A2( u2_u13_u7_n98 ) );
  NAND2_X1 u2_u13_u7_U52 (.A2( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n147 ) , .A1( u2_u13_u7_n93 ) );
  NAND2_X1 u2_u13_u7_U53 (.A1( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n127 ) , .A2( u2_u13_u7_n99 ) );
  OR2_X1 u2_u13_u7_U54 (.ZN( u2_u13_u7_n126 ) , .A2( u2_u13_u7_n152 ) , .A1( u2_u13_u7_n156 ) );
  NAND2_X1 u2_u13_u7_U55 (.A2( u2_u13_u7_n102 ) , .A1( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n133 ) );
  NAND2_X1 u2_u13_u7_U56 (.ZN( u2_u13_u7_n112 ) , .A2( u2_u13_u7_n96 ) , .A1( u2_u13_u7_n99 ) );
  NAND2_X1 u2_u13_u7_U57 (.A2( u2_u13_u7_n102 ) , .ZN( u2_u13_u7_n128 ) , .A1( u2_u13_u7_n98 ) );
  NAND2_X1 u2_u13_u7_U58 (.A1( u2_u13_u7_n100 ) , .ZN( u2_u13_u7_n113 ) , .A2( u2_u13_u7_n93 ) );
  NAND2_X1 u2_u13_u7_U59 (.A2( u2_u13_u7_n102 ) , .ZN( u2_u13_u7_n124 ) , .A1( u2_u13_u7_n96 ) );
  INV_X1 u2_u13_u7_U6 (.A( u2_u13_u7_n154 ) , .ZN( u2_u13_u7_n178 ) );
  NAND2_X1 u2_u13_u7_U60 (.ZN( u2_u13_u7_n110 ) , .A1( u2_u13_u7_n95 ) , .A2( u2_u13_u7_n96 ) );
  INV_X1 u2_u13_u7_U61 (.A( u2_u13_u7_n150 ) , .ZN( u2_u13_u7_n164 ) );
  AND2_X1 u2_u13_u7_U62 (.ZN( u2_u13_u7_n134 ) , .A1( u2_u13_u7_n93 ) , .A2( u2_u13_u7_n98 ) );
  NAND2_X1 u2_u13_u7_U63 (.A1( u2_u13_u7_n100 ) , .A2( u2_u13_u7_n102 ) , .ZN( u2_u13_u7_n129 ) );
  NAND2_X1 u2_u13_u7_U64 (.A2( u2_u13_u7_n103 ) , .ZN( u2_u13_u7_n131 ) , .A1( u2_u13_u7_n95 ) );
  NAND2_X1 u2_u13_u7_U65 (.A1( u2_u13_u7_n100 ) , .ZN( u2_u13_u7_n138 ) , .A2( u2_u13_u7_n99 ) );
  NAND2_X1 u2_u13_u7_U66 (.ZN( u2_u13_u7_n132 ) , .A1( u2_u13_u7_n93 ) , .A2( u2_u13_u7_n96 ) );
  NAND2_X1 u2_u13_u7_U67 (.A1( u2_u13_u7_n100 ) , .ZN( u2_u13_u7_n148 ) , .A2( u2_u13_u7_n95 ) );
  NOR2_X1 u2_u13_u7_U68 (.A2( u2_u13_X_47 ) , .ZN( u2_u13_u7_n150 ) , .A1( u2_u13_u7_n163 ) );
  NOR2_X1 u2_u13_u7_U69 (.A2( u2_u13_X_43 ) , .A1( u2_u13_X_44 ) , .ZN( u2_u13_u7_n103 ) );
  AOI211_X1 u2_u13_u7_U7 (.ZN( u2_u13_u7_n116 ) , .A( u2_u13_u7_n155 ) , .C1( u2_u13_u7_n161 ) , .C2( u2_u13_u7_n171 ) , .B( u2_u13_u7_n94 ) );
  NOR2_X1 u2_u13_u7_U70 (.A2( u2_u13_X_48 ) , .A1( u2_u13_u7_n166 ) , .ZN( u2_u13_u7_n95 ) );
  NOR2_X1 u2_u13_u7_U71 (.A2( u2_u13_X_45 ) , .A1( u2_u13_X_48 ) , .ZN( u2_u13_u7_n99 ) );
  NOR2_X1 u2_u13_u7_U72 (.A2( u2_u13_X_44 ) , .A1( u2_u13_u7_n167 ) , .ZN( u2_u13_u7_n98 ) );
  NOR2_X1 u2_u13_u7_U73 (.A2( u2_u13_X_46 ) , .A1( u2_u13_X_47 ) , .ZN( u2_u13_u7_n152 ) );
  AND2_X1 u2_u13_u7_U74 (.A1( u2_u13_X_47 ) , .ZN( u2_u13_u7_n156 ) , .A2( u2_u13_u7_n163 ) );
  NAND2_X1 u2_u13_u7_U75 (.A2( u2_u13_X_46 ) , .A1( u2_u13_X_47 ) , .ZN( u2_u13_u7_n125 ) );
  AND2_X1 u2_u13_u7_U76 (.A2( u2_u13_X_45 ) , .A1( u2_u13_X_48 ) , .ZN( u2_u13_u7_n102 ) );
  AND2_X1 u2_u13_u7_U77 (.A2( u2_u13_X_43 ) , .A1( u2_u13_X_44 ) , .ZN( u2_u13_u7_n96 ) );
  AND2_X1 u2_u13_u7_U78 (.A1( u2_u13_X_44 ) , .ZN( u2_u13_u7_n100 ) , .A2( u2_u13_u7_n167 ) );
  AND2_X1 u2_u13_u7_U79 (.A1( u2_u13_X_48 ) , .A2( u2_u13_u7_n166 ) , .ZN( u2_u13_u7_n93 ) );
  OAI222_X1 u2_u13_u7_U8 (.C2( u2_u13_u7_n101 ) , .B2( u2_u13_u7_n111 ) , .A1( u2_u13_u7_n113 ) , .C1( u2_u13_u7_n146 ) , .A2( u2_u13_u7_n162 ) , .B1( u2_u13_u7_n164 ) , .ZN( u2_u13_u7_n94 ) );
  INV_X1 u2_u13_u7_U80 (.A( u2_u13_X_46 ) , .ZN( u2_u13_u7_n163 ) );
  INV_X1 u2_u13_u7_U81 (.A( u2_u13_X_43 ) , .ZN( u2_u13_u7_n167 ) );
  INV_X1 u2_u13_u7_U82 (.A( u2_u13_X_45 ) , .ZN( u2_u13_u7_n166 ) );
  NAND4_X1 u2_u13_u7_U83 (.ZN( u2_out13_27 ) , .A4( u2_u13_u7_n118 ) , .A3( u2_u13_u7_n119 ) , .A2( u2_u13_u7_n120 ) , .A1( u2_u13_u7_n121 ) );
  OAI21_X1 u2_u13_u7_U84 (.ZN( u2_u13_u7_n121 ) , .B2( u2_u13_u7_n145 ) , .A( u2_u13_u7_n150 ) , .B1( u2_u13_u7_n174 ) );
  OAI21_X1 u2_u13_u7_U85 (.ZN( u2_u13_u7_n120 ) , .A( u2_u13_u7_n161 ) , .B2( u2_u13_u7_n170 ) , .B1( u2_u13_u7_n179 ) );
  NAND4_X1 u2_u13_u7_U86 (.ZN( u2_out13_21 ) , .A4( u2_u13_u7_n157 ) , .A3( u2_u13_u7_n158 ) , .A2( u2_u13_u7_n159 ) , .A1( u2_u13_u7_n160 ) );
  OAI21_X1 u2_u13_u7_U87 (.B1( u2_u13_u7_n145 ) , .ZN( u2_u13_u7_n160 ) , .A( u2_u13_u7_n161 ) , .B2( u2_u13_u7_n177 ) );
  AOI22_X1 u2_u13_u7_U88 (.B2( u2_u13_u7_n149 ) , .B1( u2_u13_u7_n150 ) , .A2( u2_u13_u7_n151 ) , .A1( u2_u13_u7_n152 ) , .ZN( u2_u13_u7_n158 ) );
  NAND4_X1 u2_u13_u7_U89 (.ZN( u2_out13_15 ) , .A4( u2_u13_u7_n142 ) , .A3( u2_u13_u7_n143 ) , .A2( u2_u13_u7_n144 ) , .A1( u2_u13_u7_n178 ) );
  OAI221_X1 u2_u13_u7_U9 (.C1( u2_u13_u7_n101 ) , .C2( u2_u13_u7_n147 ) , .ZN( u2_u13_u7_n155 ) , .B2( u2_u13_u7_n162 ) , .A( u2_u13_u7_n91 ) , .B1( u2_u13_u7_n92 ) );
  OR2_X1 u2_u13_u7_U90 (.A2( u2_u13_u7_n125 ) , .A1( u2_u13_u7_n129 ) , .ZN( u2_u13_u7_n144 ) );
  AOI22_X1 u2_u13_u7_U91 (.A2( u2_u13_u7_n126 ) , .ZN( u2_u13_u7_n143 ) , .B2( u2_u13_u7_n165 ) , .B1( u2_u13_u7_n173 ) , .A1( u2_u13_u7_n174 ) );
  NAND4_X1 u2_u13_u7_U92 (.ZN( u2_out13_5 ) , .A4( u2_u13_u7_n108 ) , .A3( u2_u13_u7_n109 ) , .A1( u2_u13_u7_n116 ) , .A2( u2_u13_u7_n123 ) );
  AOI22_X1 u2_u13_u7_U93 (.ZN( u2_u13_u7_n109 ) , .A2( u2_u13_u7_n126 ) , .B2( u2_u13_u7_n145 ) , .B1( u2_u13_u7_n156 ) , .A1( u2_u13_u7_n171 ) );
  NOR4_X1 u2_u13_u7_U94 (.A4( u2_u13_u7_n104 ) , .A3( u2_u13_u7_n105 ) , .A2( u2_u13_u7_n106 ) , .A1( u2_u13_u7_n107 ) , .ZN( u2_u13_u7_n108 ) );
  NAND3_X1 u2_u13_u7_U95 (.A3( u2_u13_u7_n146 ) , .A2( u2_u13_u7_n147 ) , .A1( u2_u13_u7_n148 ) , .ZN( u2_u13_u7_n151 ) );
  NAND3_X1 u2_u13_u7_U96 (.A3( u2_u13_u7_n131 ) , .A2( u2_u13_u7_n132 ) , .A1( u2_u13_u7_n133 ) , .ZN( u2_u13_u7_n135 ) );
  XOR2_X1 u2_u1_U13 (.B( u2_K2_42 ) , .A( u2_R0_29 ) , .Z( u2_u1_X_42 ) );
  XOR2_X1 u2_u1_U14 (.B( u2_K2_41 ) , .A( u2_R0_28 ) , .Z( u2_u1_X_41 ) );
  XOR2_X1 u2_u1_U15 (.B( u2_K2_40 ) , .A( u2_R0_27 ) , .Z( u2_u1_X_40 ) );
  XOR2_X1 u2_u1_U17 (.B( u2_K2_39 ) , .A( u2_R0_26 ) , .Z( u2_u1_X_39 ) );
  XOR2_X1 u2_u1_U18 (.B( u2_K2_38 ) , .A( u2_R0_25 ) , .Z( u2_u1_X_38 ) );
  XOR2_X1 u2_u1_U19 (.B( u2_K2_37 ) , .A( u2_R0_24 ) , .Z( u2_u1_X_37 ) );
  XOR2_X1 u2_u1_U20 (.B( u2_K2_36 ) , .A( u2_R0_25 ) , .Z( u2_u1_X_36 ) );
  XOR2_X1 u2_u1_U21 (.B( u2_K2_35 ) , .A( u2_R0_24 ) , .Z( u2_u1_X_35 ) );
  XOR2_X1 u2_u1_U22 (.B( u2_K2_34 ) , .A( u2_R0_23 ) , .Z( u2_u1_X_34 ) );
  XOR2_X1 u2_u1_U23 (.B( u2_K2_33 ) , .A( u2_R0_22 ) , .Z( u2_u1_X_33 ) );
  XOR2_X1 u2_u1_U24 (.B( u2_K2_32 ) , .A( u2_R0_21 ) , .Z( u2_u1_X_32 ) );
  XOR2_X1 u2_u1_U25 (.B( u2_K2_31 ) , .A( u2_R0_20 ) , .Z( u2_u1_X_31 ) );
  INV_X1 u2_u1_u5_U10 (.A( u2_u1_u5_n121 ) , .ZN( u2_u1_u5_n177 ) );
  NOR3_X1 u2_u1_u5_U100 (.A3( u2_u1_u5_n141 ) , .A1( u2_u1_u5_n142 ) , .ZN( u2_u1_u5_n143 ) , .A2( u2_u1_u5_n191 ) );
  NAND4_X1 u2_u1_u5_U101 (.ZN( u2_out1_4 ) , .A4( u2_u1_u5_n112 ) , .A2( u2_u1_u5_n113 ) , .A1( u2_u1_u5_n114 ) , .A3( u2_u1_u5_n195 ) );
  AOI211_X1 u2_u1_u5_U102 (.A( u2_u1_u5_n110 ) , .C1( u2_u1_u5_n111 ) , .ZN( u2_u1_u5_n112 ) , .B( u2_u1_u5_n118 ) , .C2( u2_u1_u5_n177 ) );
  AOI222_X1 u2_u1_u5_U103 (.ZN( u2_u1_u5_n113 ) , .A1( u2_u1_u5_n131 ) , .C1( u2_u1_u5_n148 ) , .B2( u2_u1_u5_n174 ) , .C2( u2_u1_u5_n178 ) , .A2( u2_u1_u5_n179 ) , .B1( u2_u1_u5_n99 ) );
  NAND3_X1 u2_u1_u5_U104 (.A2( u2_u1_u5_n154 ) , .A3( u2_u1_u5_n158 ) , .A1( u2_u1_u5_n161 ) , .ZN( u2_u1_u5_n99 ) );
  NOR2_X1 u2_u1_u5_U11 (.ZN( u2_u1_u5_n160 ) , .A2( u2_u1_u5_n173 ) , .A1( u2_u1_u5_n177 ) );
  INV_X1 u2_u1_u5_U12 (.A( u2_u1_u5_n150 ) , .ZN( u2_u1_u5_n174 ) );
  AOI21_X1 u2_u1_u5_U13 (.A( u2_u1_u5_n160 ) , .B2( u2_u1_u5_n161 ) , .ZN( u2_u1_u5_n162 ) , .B1( u2_u1_u5_n192 ) );
  INV_X1 u2_u1_u5_U14 (.A( u2_u1_u5_n159 ) , .ZN( u2_u1_u5_n192 ) );
  AOI21_X1 u2_u1_u5_U15 (.A( u2_u1_u5_n156 ) , .B2( u2_u1_u5_n157 ) , .B1( u2_u1_u5_n158 ) , .ZN( u2_u1_u5_n163 ) );
  AOI21_X1 u2_u1_u5_U16 (.B2( u2_u1_u5_n139 ) , .B1( u2_u1_u5_n140 ) , .ZN( u2_u1_u5_n141 ) , .A( u2_u1_u5_n150 ) );
  OAI21_X1 u2_u1_u5_U17 (.A( u2_u1_u5_n133 ) , .B2( u2_u1_u5_n134 ) , .B1( u2_u1_u5_n135 ) , .ZN( u2_u1_u5_n142 ) );
  OAI21_X1 u2_u1_u5_U18 (.ZN( u2_u1_u5_n133 ) , .B2( u2_u1_u5_n147 ) , .A( u2_u1_u5_n173 ) , .B1( u2_u1_u5_n188 ) );
  NAND2_X1 u2_u1_u5_U19 (.A2( u2_u1_u5_n119 ) , .A1( u2_u1_u5_n123 ) , .ZN( u2_u1_u5_n137 ) );
  INV_X1 u2_u1_u5_U20 (.A( u2_u1_u5_n155 ) , .ZN( u2_u1_u5_n194 ) );
  NAND2_X1 u2_u1_u5_U21 (.A1( u2_u1_u5_n121 ) , .ZN( u2_u1_u5_n132 ) , .A2( u2_u1_u5_n172 ) );
  NAND2_X1 u2_u1_u5_U22 (.A2( u2_u1_u5_n122 ) , .ZN( u2_u1_u5_n136 ) , .A1( u2_u1_u5_n154 ) );
  NAND2_X1 u2_u1_u5_U23 (.A2( u2_u1_u5_n119 ) , .A1( u2_u1_u5_n120 ) , .ZN( u2_u1_u5_n159 ) );
  INV_X1 u2_u1_u5_U24 (.A( u2_u1_u5_n156 ) , .ZN( u2_u1_u5_n175 ) );
  INV_X1 u2_u1_u5_U25 (.A( u2_u1_u5_n158 ) , .ZN( u2_u1_u5_n188 ) );
  INV_X1 u2_u1_u5_U26 (.A( u2_u1_u5_n152 ) , .ZN( u2_u1_u5_n179 ) );
  INV_X1 u2_u1_u5_U27 (.A( u2_u1_u5_n140 ) , .ZN( u2_u1_u5_n182 ) );
  INV_X1 u2_u1_u5_U28 (.A( u2_u1_u5_n151 ) , .ZN( u2_u1_u5_n183 ) );
  INV_X1 u2_u1_u5_U29 (.A( u2_u1_u5_n123 ) , .ZN( u2_u1_u5_n185 ) );
  NOR2_X1 u2_u1_u5_U3 (.ZN( u2_u1_u5_n134 ) , .A1( u2_u1_u5_n183 ) , .A2( u2_u1_u5_n190 ) );
  INV_X1 u2_u1_u5_U30 (.A( u2_u1_u5_n161 ) , .ZN( u2_u1_u5_n184 ) );
  INV_X1 u2_u1_u5_U31 (.A( u2_u1_u5_n139 ) , .ZN( u2_u1_u5_n189 ) );
  INV_X1 u2_u1_u5_U32 (.A( u2_u1_u5_n157 ) , .ZN( u2_u1_u5_n190 ) );
  INV_X1 u2_u1_u5_U33 (.A( u2_u1_u5_n120 ) , .ZN( u2_u1_u5_n193 ) );
  NAND2_X1 u2_u1_u5_U34 (.ZN( u2_u1_u5_n111 ) , .A1( u2_u1_u5_n140 ) , .A2( u2_u1_u5_n155 ) );
  INV_X1 u2_u1_u5_U35 (.A( u2_u1_u5_n117 ) , .ZN( u2_u1_u5_n196 ) );
  OAI221_X1 u2_u1_u5_U36 (.A( u2_u1_u5_n116 ) , .ZN( u2_u1_u5_n117 ) , .B2( u2_u1_u5_n119 ) , .C1( u2_u1_u5_n153 ) , .C2( u2_u1_u5_n158 ) , .B1( u2_u1_u5_n172 ) );
  AOI222_X1 u2_u1_u5_U37 (.ZN( u2_u1_u5_n116 ) , .B2( u2_u1_u5_n145 ) , .C1( u2_u1_u5_n148 ) , .A2( u2_u1_u5_n174 ) , .C2( u2_u1_u5_n177 ) , .B1( u2_u1_u5_n187 ) , .A1( u2_u1_u5_n193 ) );
  INV_X1 u2_u1_u5_U38 (.A( u2_u1_u5_n115 ) , .ZN( u2_u1_u5_n187 ) );
  NOR2_X1 u2_u1_u5_U39 (.ZN( u2_u1_u5_n100 ) , .A1( u2_u1_u5_n170 ) , .A2( u2_u1_u5_n180 ) );
  INV_X1 u2_u1_u5_U4 (.A( u2_u1_u5_n138 ) , .ZN( u2_u1_u5_n191 ) );
  AOI22_X1 u2_u1_u5_U40 (.B2( u2_u1_u5_n131 ) , .A2( u2_u1_u5_n146 ) , .ZN( u2_u1_u5_n169 ) , .B1( u2_u1_u5_n174 ) , .A1( u2_u1_u5_n185 ) );
  NOR2_X1 u2_u1_u5_U41 (.A1( u2_u1_u5_n146 ) , .ZN( u2_u1_u5_n150 ) , .A2( u2_u1_u5_n173 ) );
  AOI21_X1 u2_u1_u5_U42 (.A( u2_u1_u5_n118 ) , .B2( u2_u1_u5_n145 ) , .ZN( u2_u1_u5_n168 ) , .B1( u2_u1_u5_n186 ) );
  INV_X1 u2_u1_u5_U43 (.A( u2_u1_u5_n122 ) , .ZN( u2_u1_u5_n186 ) );
  NOR2_X1 u2_u1_u5_U44 (.A1( u2_u1_u5_n146 ) , .ZN( u2_u1_u5_n152 ) , .A2( u2_u1_u5_n176 ) );
  NOR2_X1 u2_u1_u5_U45 (.A1( u2_u1_u5_n115 ) , .ZN( u2_u1_u5_n118 ) , .A2( u2_u1_u5_n153 ) );
  NOR2_X1 u2_u1_u5_U46 (.A2( u2_u1_u5_n145 ) , .ZN( u2_u1_u5_n156 ) , .A1( u2_u1_u5_n174 ) );
  NOR2_X1 u2_u1_u5_U47 (.ZN( u2_u1_u5_n121 ) , .A2( u2_u1_u5_n145 ) , .A1( u2_u1_u5_n176 ) );
  AOI22_X1 u2_u1_u5_U48 (.ZN( u2_u1_u5_n114 ) , .A2( u2_u1_u5_n137 ) , .A1( u2_u1_u5_n145 ) , .B2( u2_u1_u5_n175 ) , .B1( u2_u1_u5_n193 ) );
  OAI211_X1 u2_u1_u5_U49 (.B( u2_u1_u5_n124 ) , .A( u2_u1_u5_n125 ) , .C2( u2_u1_u5_n126 ) , .C1( u2_u1_u5_n127 ) , .ZN( u2_u1_u5_n128 ) );
  OAI21_X1 u2_u1_u5_U5 (.B2( u2_u1_u5_n136 ) , .B1( u2_u1_u5_n137 ) , .ZN( u2_u1_u5_n138 ) , .A( u2_u1_u5_n177 ) );
  OAI21_X1 u2_u1_u5_U50 (.ZN( u2_u1_u5_n124 ) , .A( u2_u1_u5_n177 ) , .B2( u2_u1_u5_n183 ) , .B1( u2_u1_u5_n189 ) );
  NOR3_X1 u2_u1_u5_U51 (.ZN( u2_u1_u5_n127 ) , .A1( u2_u1_u5_n136 ) , .A3( u2_u1_u5_n148 ) , .A2( u2_u1_u5_n182 ) );
  OAI21_X1 u2_u1_u5_U52 (.ZN( u2_u1_u5_n125 ) , .A( u2_u1_u5_n174 ) , .B2( u2_u1_u5_n185 ) , .B1( u2_u1_u5_n190 ) );
  AOI21_X1 u2_u1_u5_U53 (.A( u2_u1_u5_n153 ) , .B2( u2_u1_u5_n154 ) , .B1( u2_u1_u5_n155 ) , .ZN( u2_u1_u5_n164 ) );
  AOI21_X1 u2_u1_u5_U54 (.ZN( u2_u1_u5_n110 ) , .B1( u2_u1_u5_n122 ) , .B2( u2_u1_u5_n139 ) , .A( u2_u1_u5_n153 ) );
  INV_X1 u2_u1_u5_U55 (.A( u2_u1_u5_n153 ) , .ZN( u2_u1_u5_n176 ) );
  INV_X1 u2_u1_u5_U56 (.A( u2_u1_u5_n126 ) , .ZN( u2_u1_u5_n173 ) );
  AND2_X1 u2_u1_u5_U57 (.A2( u2_u1_u5_n104 ) , .A1( u2_u1_u5_n107 ) , .ZN( u2_u1_u5_n147 ) );
  AND2_X1 u2_u1_u5_U58 (.A2( u2_u1_u5_n104 ) , .A1( u2_u1_u5_n108 ) , .ZN( u2_u1_u5_n148 ) );
  NAND2_X1 u2_u1_u5_U59 (.A1( u2_u1_u5_n105 ) , .A2( u2_u1_u5_n106 ) , .ZN( u2_u1_u5_n158 ) );
  INV_X1 u2_u1_u5_U6 (.A( u2_u1_u5_n135 ) , .ZN( u2_u1_u5_n178 ) );
  NAND2_X1 u2_u1_u5_U60 (.A2( u2_u1_u5_n108 ) , .A1( u2_u1_u5_n109 ) , .ZN( u2_u1_u5_n139 ) );
  NAND2_X1 u2_u1_u5_U61 (.A1( u2_u1_u5_n106 ) , .A2( u2_u1_u5_n108 ) , .ZN( u2_u1_u5_n119 ) );
  NAND2_X1 u2_u1_u5_U62 (.A2( u2_u1_u5_n103 ) , .A1( u2_u1_u5_n105 ) , .ZN( u2_u1_u5_n140 ) );
  NAND2_X1 u2_u1_u5_U63 (.A2( u2_u1_u5_n104 ) , .A1( u2_u1_u5_n105 ) , .ZN( u2_u1_u5_n155 ) );
  NAND2_X1 u2_u1_u5_U64 (.A2( u2_u1_u5_n106 ) , .A1( u2_u1_u5_n107 ) , .ZN( u2_u1_u5_n122 ) );
  NAND2_X1 u2_u1_u5_U65 (.A2( u2_u1_u5_n100 ) , .A1( u2_u1_u5_n106 ) , .ZN( u2_u1_u5_n115 ) );
  NAND2_X1 u2_u1_u5_U66 (.A2( u2_u1_u5_n100 ) , .A1( u2_u1_u5_n103 ) , .ZN( u2_u1_u5_n161 ) );
  NAND2_X1 u2_u1_u5_U67 (.A1( u2_u1_u5_n105 ) , .A2( u2_u1_u5_n109 ) , .ZN( u2_u1_u5_n154 ) );
  INV_X1 u2_u1_u5_U68 (.A( u2_u1_u5_n146 ) , .ZN( u2_u1_u5_n172 ) );
  NAND2_X1 u2_u1_u5_U69 (.A1( u2_u1_u5_n103 ) , .A2( u2_u1_u5_n108 ) , .ZN( u2_u1_u5_n123 ) );
  OAI22_X1 u2_u1_u5_U7 (.B2( u2_u1_u5_n149 ) , .B1( u2_u1_u5_n150 ) , .A2( u2_u1_u5_n151 ) , .A1( u2_u1_u5_n152 ) , .ZN( u2_u1_u5_n165 ) );
  NAND2_X1 u2_u1_u5_U70 (.A2( u2_u1_u5_n103 ) , .A1( u2_u1_u5_n107 ) , .ZN( u2_u1_u5_n151 ) );
  NAND2_X1 u2_u1_u5_U71 (.A2( u2_u1_u5_n107 ) , .A1( u2_u1_u5_n109 ) , .ZN( u2_u1_u5_n120 ) );
  NAND2_X1 u2_u1_u5_U72 (.A2( u2_u1_u5_n100 ) , .A1( u2_u1_u5_n109 ) , .ZN( u2_u1_u5_n157 ) );
  AND2_X1 u2_u1_u5_U73 (.A2( u2_u1_u5_n100 ) , .A1( u2_u1_u5_n104 ) , .ZN( u2_u1_u5_n131 ) );
  INV_X1 u2_u1_u5_U74 (.A( u2_u1_u5_n102 ) , .ZN( u2_u1_u5_n195 ) );
  OAI221_X1 u2_u1_u5_U75 (.A( u2_u1_u5_n101 ) , .ZN( u2_u1_u5_n102 ) , .C2( u2_u1_u5_n115 ) , .C1( u2_u1_u5_n126 ) , .B1( u2_u1_u5_n134 ) , .B2( u2_u1_u5_n160 ) );
  OAI21_X1 u2_u1_u5_U76 (.ZN( u2_u1_u5_n101 ) , .B1( u2_u1_u5_n137 ) , .A( u2_u1_u5_n146 ) , .B2( u2_u1_u5_n147 ) );
  NOR2_X1 u2_u1_u5_U77 (.A2( u2_u1_X_34 ) , .A1( u2_u1_X_35 ) , .ZN( u2_u1_u5_n145 ) );
  NOR2_X1 u2_u1_u5_U78 (.A2( u2_u1_X_34 ) , .ZN( u2_u1_u5_n146 ) , .A1( u2_u1_u5_n171 ) );
  NOR2_X1 u2_u1_u5_U79 (.A2( u2_u1_X_31 ) , .A1( u2_u1_X_32 ) , .ZN( u2_u1_u5_n103 ) );
  NOR3_X1 u2_u1_u5_U8 (.A2( u2_u1_u5_n147 ) , .A1( u2_u1_u5_n148 ) , .ZN( u2_u1_u5_n149 ) , .A3( u2_u1_u5_n194 ) );
  NOR2_X1 u2_u1_u5_U80 (.A2( u2_u1_X_36 ) , .ZN( u2_u1_u5_n105 ) , .A1( u2_u1_u5_n180 ) );
  NOR2_X1 u2_u1_u5_U81 (.A2( u2_u1_X_33 ) , .ZN( u2_u1_u5_n108 ) , .A1( u2_u1_u5_n170 ) );
  NOR2_X1 u2_u1_u5_U82 (.A2( u2_u1_X_33 ) , .A1( u2_u1_X_36 ) , .ZN( u2_u1_u5_n107 ) );
  NOR2_X1 u2_u1_u5_U83 (.A2( u2_u1_X_31 ) , .ZN( u2_u1_u5_n104 ) , .A1( u2_u1_u5_n181 ) );
  NAND2_X1 u2_u1_u5_U84 (.A2( u2_u1_X_34 ) , .A1( u2_u1_X_35 ) , .ZN( u2_u1_u5_n153 ) );
  NAND2_X1 u2_u1_u5_U85 (.A1( u2_u1_X_34 ) , .ZN( u2_u1_u5_n126 ) , .A2( u2_u1_u5_n171 ) );
  AND2_X1 u2_u1_u5_U86 (.A1( u2_u1_X_31 ) , .A2( u2_u1_X_32 ) , .ZN( u2_u1_u5_n106 ) );
  AND2_X1 u2_u1_u5_U87 (.A1( u2_u1_X_31 ) , .ZN( u2_u1_u5_n109 ) , .A2( u2_u1_u5_n181 ) );
  INV_X1 u2_u1_u5_U88 (.A( u2_u1_X_33 ) , .ZN( u2_u1_u5_n180 ) );
  INV_X1 u2_u1_u5_U89 (.A( u2_u1_X_35 ) , .ZN( u2_u1_u5_n171 ) );
  NOR2_X1 u2_u1_u5_U9 (.ZN( u2_u1_u5_n135 ) , .A1( u2_u1_u5_n173 ) , .A2( u2_u1_u5_n176 ) );
  INV_X1 u2_u1_u5_U90 (.A( u2_u1_X_36 ) , .ZN( u2_u1_u5_n170 ) );
  INV_X1 u2_u1_u5_U91 (.A( u2_u1_X_32 ) , .ZN( u2_u1_u5_n181 ) );
  NAND4_X1 u2_u1_u5_U92 (.ZN( u2_out1_29 ) , .A4( u2_u1_u5_n129 ) , .A3( u2_u1_u5_n130 ) , .A2( u2_u1_u5_n168 ) , .A1( u2_u1_u5_n196 ) );
  AOI221_X1 u2_u1_u5_U93 (.A( u2_u1_u5_n128 ) , .ZN( u2_u1_u5_n129 ) , .C2( u2_u1_u5_n132 ) , .B2( u2_u1_u5_n159 ) , .B1( u2_u1_u5_n176 ) , .C1( u2_u1_u5_n184 ) );
  AOI222_X1 u2_u1_u5_U94 (.ZN( u2_u1_u5_n130 ) , .A2( u2_u1_u5_n146 ) , .B1( u2_u1_u5_n147 ) , .C2( u2_u1_u5_n175 ) , .B2( u2_u1_u5_n179 ) , .A1( u2_u1_u5_n188 ) , .C1( u2_u1_u5_n194 ) );
  NAND4_X1 u2_u1_u5_U95 (.ZN( u2_out1_19 ) , .A4( u2_u1_u5_n166 ) , .A3( u2_u1_u5_n167 ) , .A2( u2_u1_u5_n168 ) , .A1( u2_u1_u5_n169 ) );
  AOI22_X1 u2_u1_u5_U96 (.B2( u2_u1_u5_n145 ) , .A2( u2_u1_u5_n146 ) , .ZN( u2_u1_u5_n167 ) , .B1( u2_u1_u5_n182 ) , .A1( u2_u1_u5_n189 ) );
  NOR4_X1 u2_u1_u5_U97 (.A4( u2_u1_u5_n162 ) , .A3( u2_u1_u5_n163 ) , .A2( u2_u1_u5_n164 ) , .A1( u2_u1_u5_n165 ) , .ZN( u2_u1_u5_n166 ) );
  NAND4_X1 u2_u1_u5_U98 (.ZN( u2_out1_11 ) , .A4( u2_u1_u5_n143 ) , .A3( u2_u1_u5_n144 ) , .A2( u2_u1_u5_n169 ) , .A1( u2_u1_u5_n196 ) );
  AOI22_X1 u2_u1_u5_U99 (.A2( u2_u1_u5_n132 ) , .ZN( u2_u1_u5_n144 ) , .B2( u2_u1_u5_n145 ) , .B1( u2_u1_u5_n184 ) , .A1( u2_u1_u5_n194 ) );
  AOI22_X1 u2_u1_u6_U10 (.A2( u2_u1_u6_n151 ) , .B2( u2_u1_u6_n161 ) , .A1( u2_u1_u6_n167 ) , .B1( u2_u1_u6_n170 ) , .ZN( u2_u1_u6_n89 ) );
  AOI21_X1 u2_u1_u6_U11 (.B1( u2_u1_u6_n107 ) , .B2( u2_u1_u6_n132 ) , .A( u2_u1_u6_n158 ) , .ZN( u2_u1_u6_n88 ) );
  AOI21_X1 u2_u1_u6_U12 (.B2( u2_u1_u6_n147 ) , .B1( u2_u1_u6_n148 ) , .ZN( u2_u1_u6_n149 ) , .A( u2_u1_u6_n158 ) );
  AOI21_X1 u2_u1_u6_U13 (.ZN( u2_u1_u6_n106 ) , .A( u2_u1_u6_n142 ) , .B2( u2_u1_u6_n159 ) , .B1( u2_u1_u6_n164 ) );
  INV_X1 u2_u1_u6_U14 (.A( u2_u1_u6_n155 ) , .ZN( u2_u1_u6_n161 ) );
  INV_X1 u2_u1_u6_U15 (.A( u2_u1_u6_n128 ) , .ZN( u2_u1_u6_n164 ) );
  NAND2_X1 u2_u1_u6_U16 (.ZN( u2_u1_u6_n110 ) , .A1( u2_u1_u6_n122 ) , .A2( u2_u1_u6_n129 ) );
  NAND2_X1 u2_u1_u6_U17 (.ZN( u2_u1_u6_n124 ) , .A2( u2_u1_u6_n146 ) , .A1( u2_u1_u6_n148 ) );
  INV_X1 u2_u1_u6_U18 (.A( u2_u1_u6_n132 ) , .ZN( u2_u1_u6_n171 ) );
  AND2_X1 u2_u1_u6_U19 (.A1( u2_u1_u6_n100 ) , .ZN( u2_u1_u6_n130 ) , .A2( u2_u1_u6_n147 ) );
  INV_X1 u2_u1_u6_U20 (.A( u2_u1_u6_n127 ) , .ZN( u2_u1_u6_n173 ) );
  INV_X1 u2_u1_u6_U21 (.A( u2_u1_u6_n121 ) , .ZN( u2_u1_u6_n167 ) );
  INV_X1 u2_u1_u6_U22 (.A( u2_u1_u6_n100 ) , .ZN( u2_u1_u6_n169 ) );
  INV_X1 u2_u1_u6_U23 (.A( u2_u1_u6_n123 ) , .ZN( u2_u1_u6_n170 ) );
  INV_X1 u2_u1_u6_U24 (.A( u2_u1_u6_n113 ) , .ZN( u2_u1_u6_n168 ) );
  AND2_X1 u2_u1_u6_U25 (.A1( u2_u1_u6_n107 ) , .A2( u2_u1_u6_n119 ) , .ZN( u2_u1_u6_n133 ) );
  AND2_X1 u2_u1_u6_U26 (.A2( u2_u1_u6_n121 ) , .A1( u2_u1_u6_n122 ) , .ZN( u2_u1_u6_n131 ) );
  AND3_X1 u2_u1_u6_U27 (.ZN( u2_u1_u6_n120 ) , .A2( u2_u1_u6_n127 ) , .A1( u2_u1_u6_n132 ) , .A3( u2_u1_u6_n145 ) );
  INV_X1 u2_u1_u6_U28 (.A( u2_u1_u6_n146 ) , .ZN( u2_u1_u6_n163 ) );
  AOI222_X1 u2_u1_u6_U29 (.ZN( u2_u1_u6_n114 ) , .A1( u2_u1_u6_n118 ) , .A2( u2_u1_u6_n126 ) , .B2( u2_u1_u6_n151 ) , .C2( u2_u1_u6_n159 ) , .C1( u2_u1_u6_n168 ) , .B1( u2_u1_u6_n169 ) );
  INV_X1 u2_u1_u6_U3 (.A( u2_u1_u6_n110 ) , .ZN( u2_u1_u6_n166 ) );
  NOR2_X1 u2_u1_u6_U30 (.A1( u2_u1_u6_n162 ) , .A2( u2_u1_u6_n165 ) , .ZN( u2_u1_u6_n98 ) );
  AOI211_X1 u2_u1_u6_U31 (.B( u2_u1_u6_n134 ) , .A( u2_u1_u6_n135 ) , .C1( u2_u1_u6_n136 ) , .ZN( u2_u1_u6_n137 ) , .C2( u2_u1_u6_n151 ) );
  AOI21_X1 u2_u1_u6_U32 (.B1( u2_u1_u6_n131 ) , .ZN( u2_u1_u6_n135 ) , .A( u2_u1_u6_n144 ) , .B2( u2_u1_u6_n146 ) );
  NAND4_X1 u2_u1_u6_U33 (.A4( u2_u1_u6_n127 ) , .A3( u2_u1_u6_n128 ) , .A2( u2_u1_u6_n129 ) , .A1( u2_u1_u6_n130 ) , .ZN( u2_u1_u6_n136 ) );
  AOI21_X1 u2_u1_u6_U34 (.B2( u2_u1_u6_n132 ) , .B1( u2_u1_u6_n133 ) , .ZN( u2_u1_u6_n134 ) , .A( u2_u1_u6_n158 ) );
  NAND2_X1 u2_u1_u6_U35 (.A1( u2_u1_u6_n144 ) , .ZN( u2_u1_u6_n151 ) , .A2( u2_u1_u6_n158 ) );
  NAND2_X1 u2_u1_u6_U36 (.ZN( u2_u1_u6_n132 ) , .A1( u2_u1_u6_n91 ) , .A2( u2_u1_u6_n97 ) );
  AOI22_X1 u2_u1_u6_U37 (.B2( u2_u1_u6_n110 ) , .B1( u2_u1_u6_n111 ) , .A1( u2_u1_u6_n112 ) , .ZN( u2_u1_u6_n115 ) , .A2( u2_u1_u6_n161 ) );
  NAND4_X1 u2_u1_u6_U38 (.A3( u2_u1_u6_n109 ) , .ZN( u2_u1_u6_n112 ) , .A4( u2_u1_u6_n132 ) , .A2( u2_u1_u6_n147 ) , .A1( u2_u1_u6_n166 ) );
  NOR2_X1 u2_u1_u6_U39 (.ZN( u2_u1_u6_n109 ) , .A1( u2_u1_u6_n170 ) , .A2( u2_u1_u6_n173 ) );
  INV_X1 u2_u1_u6_U4 (.A( u2_u1_u6_n142 ) , .ZN( u2_u1_u6_n174 ) );
  NOR2_X1 u2_u1_u6_U40 (.A2( u2_u1_u6_n126 ) , .ZN( u2_u1_u6_n155 ) , .A1( u2_u1_u6_n160 ) );
  NAND2_X1 u2_u1_u6_U41 (.ZN( u2_u1_u6_n146 ) , .A2( u2_u1_u6_n94 ) , .A1( u2_u1_u6_n99 ) );
  AOI21_X1 u2_u1_u6_U42 (.A( u2_u1_u6_n144 ) , .B2( u2_u1_u6_n145 ) , .B1( u2_u1_u6_n146 ) , .ZN( u2_u1_u6_n150 ) );
  INV_X1 u2_u1_u6_U43 (.A( u2_u1_u6_n111 ) , .ZN( u2_u1_u6_n158 ) );
  NAND2_X1 u2_u1_u6_U44 (.ZN( u2_u1_u6_n127 ) , .A1( u2_u1_u6_n91 ) , .A2( u2_u1_u6_n92 ) );
  NAND2_X1 u2_u1_u6_U45 (.ZN( u2_u1_u6_n129 ) , .A2( u2_u1_u6_n95 ) , .A1( u2_u1_u6_n96 ) );
  INV_X1 u2_u1_u6_U46 (.A( u2_u1_u6_n144 ) , .ZN( u2_u1_u6_n159 ) );
  NAND2_X1 u2_u1_u6_U47 (.ZN( u2_u1_u6_n145 ) , .A2( u2_u1_u6_n97 ) , .A1( u2_u1_u6_n98 ) );
  NAND2_X1 u2_u1_u6_U48 (.ZN( u2_u1_u6_n148 ) , .A2( u2_u1_u6_n92 ) , .A1( u2_u1_u6_n94 ) );
  NAND2_X1 u2_u1_u6_U49 (.ZN( u2_u1_u6_n108 ) , .A2( u2_u1_u6_n139 ) , .A1( u2_u1_u6_n144 ) );
  NAND2_X1 u2_u1_u6_U5 (.A2( u2_u1_u6_n143 ) , .ZN( u2_u1_u6_n152 ) , .A1( u2_u1_u6_n166 ) );
  NAND2_X1 u2_u1_u6_U50 (.ZN( u2_u1_u6_n121 ) , .A2( u2_u1_u6_n95 ) , .A1( u2_u1_u6_n97 ) );
  NAND2_X1 u2_u1_u6_U51 (.ZN( u2_u1_u6_n107 ) , .A2( u2_u1_u6_n92 ) , .A1( u2_u1_u6_n95 ) );
  AND2_X1 u2_u1_u6_U52 (.ZN( u2_u1_u6_n118 ) , .A2( u2_u1_u6_n91 ) , .A1( u2_u1_u6_n99 ) );
  NAND2_X1 u2_u1_u6_U53 (.ZN( u2_u1_u6_n147 ) , .A2( u2_u1_u6_n98 ) , .A1( u2_u1_u6_n99 ) );
  NAND2_X1 u2_u1_u6_U54 (.ZN( u2_u1_u6_n128 ) , .A1( u2_u1_u6_n94 ) , .A2( u2_u1_u6_n96 ) );
  NAND2_X1 u2_u1_u6_U55 (.ZN( u2_u1_u6_n119 ) , .A2( u2_u1_u6_n95 ) , .A1( u2_u1_u6_n99 ) );
  NAND2_X1 u2_u1_u6_U56 (.ZN( u2_u1_u6_n123 ) , .A2( u2_u1_u6_n91 ) , .A1( u2_u1_u6_n96 ) );
  NAND2_X1 u2_u1_u6_U57 (.ZN( u2_u1_u6_n100 ) , .A2( u2_u1_u6_n92 ) , .A1( u2_u1_u6_n98 ) );
  NAND2_X1 u2_u1_u6_U58 (.ZN( u2_u1_u6_n122 ) , .A1( u2_u1_u6_n94 ) , .A2( u2_u1_u6_n97 ) );
  INV_X1 u2_u1_u6_U59 (.A( u2_u1_u6_n139 ) , .ZN( u2_u1_u6_n160 ) );
  AOI22_X1 u2_u1_u6_U6 (.B2( u2_u1_u6_n101 ) , .A1( u2_u1_u6_n102 ) , .ZN( u2_u1_u6_n103 ) , .B1( u2_u1_u6_n160 ) , .A2( u2_u1_u6_n161 ) );
  NAND2_X1 u2_u1_u6_U60 (.ZN( u2_u1_u6_n113 ) , .A1( u2_u1_u6_n96 ) , .A2( u2_u1_u6_n98 ) );
  NOR2_X1 u2_u1_u6_U61 (.A2( u2_u1_X_40 ) , .A1( u2_u1_X_41 ) , .ZN( u2_u1_u6_n126 ) );
  NOR2_X1 u2_u1_u6_U62 (.A2( u2_u1_X_39 ) , .A1( u2_u1_X_42 ) , .ZN( u2_u1_u6_n92 ) );
  NOR2_X1 u2_u1_u6_U63 (.A2( u2_u1_X_39 ) , .A1( u2_u1_u6_n156 ) , .ZN( u2_u1_u6_n97 ) );
  NOR2_X1 u2_u1_u6_U64 (.A2( u2_u1_X_38 ) , .A1( u2_u1_u6_n165 ) , .ZN( u2_u1_u6_n95 ) );
  NOR2_X1 u2_u1_u6_U65 (.A2( u2_u1_X_41 ) , .ZN( u2_u1_u6_n111 ) , .A1( u2_u1_u6_n157 ) );
  NOR2_X1 u2_u1_u6_U66 (.A2( u2_u1_X_37 ) , .A1( u2_u1_u6_n162 ) , .ZN( u2_u1_u6_n94 ) );
  NOR2_X1 u2_u1_u6_U67 (.A2( u2_u1_X_37 ) , .A1( u2_u1_X_38 ) , .ZN( u2_u1_u6_n91 ) );
  NAND2_X1 u2_u1_u6_U68 (.A1( u2_u1_X_41 ) , .ZN( u2_u1_u6_n144 ) , .A2( u2_u1_u6_n157 ) );
  NAND2_X1 u2_u1_u6_U69 (.A2( u2_u1_X_40 ) , .A1( u2_u1_X_41 ) , .ZN( u2_u1_u6_n139 ) );
  NOR2_X1 u2_u1_u6_U7 (.A1( u2_u1_u6_n118 ) , .ZN( u2_u1_u6_n143 ) , .A2( u2_u1_u6_n168 ) );
  AND2_X1 u2_u1_u6_U70 (.A1( u2_u1_X_39 ) , .A2( u2_u1_u6_n156 ) , .ZN( u2_u1_u6_n96 ) );
  AND2_X1 u2_u1_u6_U71 (.A1( u2_u1_X_39 ) , .A2( u2_u1_X_42 ) , .ZN( u2_u1_u6_n99 ) );
  INV_X1 u2_u1_u6_U72 (.A( u2_u1_X_40 ) , .ZN( u2_u1_u6_n157 ) );
  INV_X1 u2_u1_u6_U73 (.A( u2_u1_X_37 ) , .ZN( u2_u1_u6_n165 ) );
  INV_X1 u2_u1_u6_U74 (.A( u2_u1_X_38 ) , .ZN( u2_u1_u6_n162 ) );
  INV_X1 u2_u1_u6_U75 (.A( u2_u1_X_42 ) , .ZN( u2_u1_u6_n156 ) );
  NAND4_X1 u2_u1_u6_U76 (.ZN( u2_out1_32 ) , .A4( u2_u1_u6_n103 ) , .A3( u2_u1_u6_n104 ) , .A2( u2_u1_u6_n105 ) , .A1( u2_u1_u6_n106 ) );
  AOI22_X1 u2_u1_u6_U77 (.ZN( u2_u1_u6_n105 ) , .A2( u2_u1_u6_n108 ) , .A1( u2_u1_u6_n118 ) , .B2( u2_u1_u6_n126 ) , .B1( u2_u1_u6_n171 ) );
  AOI22_X1 u2_u1_u6_U78 (.ZN( u2_u1_u6_n104 ) , .A1( u2_u1_u6_n111 ) , .B1( u2_u1_u6_n124 ) , .B2( u2_u1_u6_n151 ) , .A2( u2_u1_u6_n93 ) );
  NAND4_X1 u2_u1_u6_U79 (.ZN( u2_out1_12 ) , .A4( u2_u1_u6_n114 ) , .A3( u2_u1_u6_n115 ) , .A2( u2_u1_u6_n116 ) , .A1( u2_u1_u6_n117 ) );
  OAI21_X1 u2_u1_u6_U8 (.A( u2_u1_u6_n159 ) , .B1( u2_u1_u6_n169 ) , .B2( u2_u1_u6_n173 ) , .ZN( u2_u1_u6_n90 ) );
  OAI22_X1 u2_u1_u6_U80 (.B2( u2_u1_u6_n111 ) , .ZN( u2_u1_u6_n116 ) , .B1( u2_u1_u6_n126 ) , .A2( u2_u1_u6_n164 ) , .A1( u2_u1_u6_n167 ) );
  OAI21_X1 u2_u1_u6_U81 (.A( u2_u1_u6_n108 ) , .ZN( u2_u1_u6_n117 ) , .B2( u2_u1_u6_n141 ) , .B1( u2_u1_u6_n163 ) );
  OAI211_X1 u2_u1_u6_U82 (.ZN( u2_out1_22 ) , .B( u2_u1_u6_n137 ) , .A( u2_u1_u6_n138 ) , .C2( u2_u1_u6_n139 ) , .C1( u2_u1_u6_n140 ) );
  AND4_X1 u2_u1_u6_U83 (.A3( u2_u1_u6_n119 ) , .A1( u2_u1_u6_n120 ) , .A4( u2_u1_u6_n129 ) , .ZN( u2_u1_u6_n140 ) , .A2( u2_u1_u6_n143 ) );
  AOI22_X1 u2_u1_u6_U84 (.B1( u2_u1_u6_n124 ) , .A2( u2_u1_u6_n125 ) , .A1( u2_u1_u6_n126 ) , .ZN( u2_u1_u6_n138 ) , .B2( u2_u1_u6_n161 ) );
  OAI211_X1 u2_u1_u6_U85 (.ZN( u2_out1_7 ) , .B( u2_u1_u6_n153 ) , .C2( u2_u1_u6_n154 ) , .C1( u2_u1_u6_n155 ) , .A( u2_u1_u6_n174 ) );
  NOR3_X1 u2_u1_u6_U86 (.A1( u2_u1_u6_n141 ) , .ZN( u2_u1_u6_n154 ) , .A3( u2_u1_u6_n164 ) , .A2( u2_u1_u6_n171 ) );
  AOI211_X1 u2_u1_u6_U87 (.B( u2_u1_u6_n149 ) , .A( u2_u1_u6_n150 ) , .C2( u2_u1_u6_n151 ) , .C1( u2_u1_u6_n152 ) , .ZN( u2_u1_u6_n153 ) );
  NAND3_X1 u2_u1_u6_U88 (.A2( u2_u1_u6_n123 ) , .ZN( u2_u1_u6_n125 ) , .A1( u2_u1_u6_n130 ) , .A3( u2_u1_u6_n131 ) );
  NAND3_X1 u2_u1_u6_U89 (.A3( u2_u1_u6_n133 ) , .ZN( u2_u1_u6_n141 ) , .A1( u2_u1_u6_n145 ) , .A2( u2_u1_u6_n148 ) );
  INV_X1 u2_u1_u6_U9 (.ZN( u2_u1_u6_n172 ) , .A( u2_u1_u6_n88 ) );
  NAND3_X1 u2_u1_u6_U90 (.ZN( u2_u1_u6_n101 ) , .A3( u2_u1_u6_n107 ) , .A2( u2_u1_u6_n121 ) , .A1( u2_u1_u6_n127 ) );
  NAND3_X1 u2_u1_u6_U91 (.ZN( u2_u1_u6_n102 ) , .A3( u2_u1_u6_n130 ) , .A2( u2_u1_u6_n145 ) , .A1( u2_u1_u6_n166 ) );
  NAND3_X1 u2_u1_u6_U92 (.A3( u2_u1_u6_n113 ) , .A1( u2_u1_u6_n119 ) , .A2( u2_u1_u6_n123 ) , .ZN( u2_u1_u6_n93 ) );
  NAND3_X1 u2_u1_u6_U93 (.ZN( u2_u1_u6_n142 ) , .A2( u2_u1_u6_n172 ) , .A3( u2_u1_u6_n89 ) , .A1( u2_u1_u6_n90 ) );
  XOR2_X1 u2_u4_U1 (.B( u2_K5_9 ) , .A( u2_R3_6 ) , .Z( u2_u4_X_9 ) );
  XOR2_X1 u2_u4_U16 (.B( u2_K5_3 ) , .A( u2_R3_2 ) , .Z( u2_u4_X_3 ) );
  XOR2_X1 u2_u4_U2 (.B( u2_K5_8 ) , .A( u2_R3_5 ) , .Z( u2_u4_X_8 ) );
  XOR2_X1 u2_u4_U26 (.B( u2_K5_30 ) , .A( u2_R3_21 ) , .Z( u2_u4_X_30 ) );
  XOR2_X1 u2_u4_U27 (.B( u2_K5_2 ) , .A( u2_R3_1 ) , .Z( u2_u4_X_2 ) );
  XOR2_X1 u2_u4_U28 (.B( u2_K5_29 ) , .A( u2_R3_20 ) , .Z( u2_u4_X_29 ) );
  XOR2_X1 u2_u4_U29 (.B( u2_K5_28 ) , .A( u2_R3_19 ) , .Z( u2_u4_X_28 ) );
  XOR2_X1 u2_u4_U3 (.B( u2_K5_7 ) , .A( u2_R3_4 ) , .Z( u2_u4_X_7 ) );
  XOR2_X1 u2_u4_U30 (.B( u2_K5_27 ) , .A( u2_R3_18 ) , .Z( u2_u4_X_27 ) );
  XOR2_X1 u2_u4_U31 (.B( u2_K5_26 ) , .A( u2_R3_17 ) , .Z( u2_u4_X_26 ) );
  XOR2_X1 u2_u4_U32 (.B( u2_K5_25 ) , .A( u2_R3_16 ) , .Z( u2_u4_X_25 ) );
  XOR2_X1 u2_u4_U33 (.B( u2_K5_24 ) , .A( u2_R3_17 ) , .Z( u2_u4_X_24 ) );
  XOR2_X1 u2_u4_U34 (.B( u2_K5_23 ) , .A( u2_R3_16 ) , .Z( u2_u4_X_23 ) );
  XOR2_X1 u2_u4_U35 (.B( u2_K5_22 ) , .A( u2_R3_15 ) , .Z( u2_u4_X_22 ) );
  XOR2_X1 u2_u4_U36 (.B( u2_K5_21 ) , .A( u2_R3_14 ) , .Z( u2_u4_X_21 ) );
  XOR2_X1 u2_u4_U37 (.B( u2_K5_20 ) , .A( u2_R3_13 ) , .Z( u2_u4_X_20 ) );
  XOR2_X1 u2_u4_U38 (.B( u2_K5_1 ) , .A( u2_R3_32 ) , .Z( u2_u4_X_1 ) );
  XOR2_X1 u2_u4_U39 (.B( u2_K5_19 ) , .A( u2_R3_12 ) , .Z( u2_u4_X_19 ) );
  XOR2_X1 u2_u4_U4 (.B( u2_K5_6 ) , .A( u2_R3_5 ) , .Z( u2_u4_X_6 ) );
  XOR2_X1 u2_u4_U40 (.B( u2_K5_18 ) , .A( u2_R3_13 ) , .Z( u2_u4_X_18 ) );
  XOR2_X1 u2_u4_U41 (.B( u2_K5_17 ) , .A( u2_R3_12 ) , .Z( u2_u4_X_17 ) );
  XOR2_X1 u2_u4_U42 (.B( u2_K5_16 ) , .A( u2_R3_11 ) , .Z( u2_u4_X_16 ) );
  XOR2_X1 u2_u4_U43 (.B( u2_K5_15 ) , .A( u2_R3_10 ) , .Z( u2_u4_X_15 ) );
  XOR2_X1 u2_u4_U44 (.B( u2_K5_14 ) , .A( u2_R3_9 ) , .Z( u2_u4_X_14 ) );
  XOR2_X1 u2_u4_U45 (.B( u2_K5_13 ) , .A( u2_R3_8 ) , .Z( u2_u4_X_13 ) );
  XOR2_X1 u2_u4_U46 (.B( u2_K5_12 ) , .A( u2_R3_9 ) , .Z( u2_u4_X_12 ) );
  XOR2_X1 u2_u4_U47 (.B( u2_K5_11 ) , .A( u2_R3_8 ) , .Z( u2_u4_X_11 ) );
  XOR2_X1 u2_u4_U48 (.B( u2_K5_10 ) , .A( u2_R3_7 ) , .Z( u2_u4_X_10 ) );
  XOR2_X1 u2_u4_U5 (.B( u2_K5_5 ) , .A( u2_R3_4 ) , .Z( u2_u4_X_5 ) );
  XOR2_X1 u2_u4_U6 (.B( u2_K5_4 ) , .A( u2_R3_3 ) , .Z( u2_u4_X_4 ) );
  AND3_X1 u2_u4_u0_U10 (.A2( u2_u4_u0_n112 ) , .ZN( u2_u4_u0_n127 ) , .A3( u2_u4_u0_n130 ) , .A1( u2_u4_u0_n148 ) );
  NAND2_X1 u2_u4_u0_U11 (.ZN( u2_u4_u0_n113 ) , .A1( u2_u4_u0_n139 ) , .A2( u2_u4_u0_n149 ) );
  AND2_X1 u2_u4_u0_U12 (.ZN( u2_u4_u0_n107 ) , .A1( u2_u4_u0_n130 ) , .A2( u2_u4_u0_n140 ) );
  AND2_X1 u2_u4_u0_U13 (.A2( u2_u4_u0_n129 ) , .A1( u2_u4_u0_n130 ) , .ZN( u2_u4_u0_n151 ) );
  AND2_X1 u2_u4_u0_U14 (.A1( u2_u4_u0_n108 ) , .A2( u2_u4_u0_n125 ) , .ZN( u2_u4_u0_n145 ) );
  INV_X1 u2_u4_u0_U15 (.A( u2_u4_u0_n143 ) , .ZN( u2_u4_u0_n173 ) );
  NOR2_X1 u2_u4_u0_U16 (.A2( u2_u4_u0_n136 ) , .ZN( u2_u4_u0_n147 ) , .A1( u2_u4_u0_n160 ) );
  NOR2_X1 u2_u4_u0_U17 (.A1( u2_u4_u0_n163 ) , .A2( u2_u4_u0_n164 ) , .ZN( u2_u4_u0_n95 ) );
  AOI21_X1 u2_u4_u0_U18 (.B1( u2_u4_u0_n103 ) , .ZN( u2_u4_u0_n132 ) , .A( u2_u4_u0_n165 ) , .B2( u2_u4_u0_n93 ) );
  INV_X1 u2_u4_u0_U19 (.A( u2_u4_u0_n142 ) , .ZN( u2_u4_u0_n165 ) );
  OAI221_X1 u2_u4_u0_U20 (.C1( u2_u4_u0_n121 ) , .ZN( u2_u4_u0_n122 ) , .B2( u2_u4_u0_n127 ) , .A( u2_u4_u0_n143 ) , .B1( u2_u4_u0_n144 ) , .C2( u2_u4_u0_n147 ) );
  OAI22_X1 u2_u4_u0_U21 (.B1( u2_u4_u0_n125 ) , .ZN( u2_u4_u0_n126 ) , .A1( u2_u4_u0_n138 ) , .A2( u2_u4_u0_n146 ) , .B2( u2_u4_u0_n147 ) );
  OAI22_X1 u2_u4_u0_U22 (.B1( u2_u4_u0_n131 ) , .A1( u2_u4_u0_n144 ) , .B2( u2_u4_u0_n147 ) , .A2( u2_u4_u0_n90 ) , .ZN( u2_u4_u0_n91 ) );
  AND3_X1 u2_u4_u0_U23 (.A3( u2_u4_u0_n121 ) , .A2( u2_u4_u0_n125 ) , .A1( u2_u4_u0_n148 ) , .ZN( u2_u4_u0_n90 ) );
  NAND2_X1 u2_u4_u0_U24 (.A1( u2_u4_u0_n100 ) , .A2( u2_u4_u0_n103 ) , .ZN( u2_u4_u0_n125 ) );
  INV_X1 u2_u4_u0_U25 (.A( u2_u4_u0_n136 ) , .ZN( u2_u4_u0_n161 ) );
  NOR2_X1 u2_u4_u0_U26 (.A1( u2_u4_u0_n120 ) , .ZN( u2_u4_u0_n143 ) , .A2( u2_u4_u0_n167 ) );
  OAI221_X1 u2_u4_u0_U27 (.C1( u2_u4_u0_n112 ) , .ZN( u2_u4_u0_n120 ) , .B1( u2_u4_u0_n138 ) , .B2( u2_u4_u0_n141 ) , .C2( u2_u4_u0_n147 ) , .A( u2_u4_u0_n172 ) );
  AOI211_X1 u2_u4_u0_U28 (.B( u2_u4_u0_n115 ) , .A( u2_u4_u0_n116 ) , .C2( u2_u4_u0_n117 ) , .C1( u2_u4_u0_n118 ) , .ZN( u2_u4_u0_n119 ) );
  AOI22_X1 u2_u4_u0_U29 (.B2( u2_u4_u0_n109 ) , .A2( u2_u4_u0_n110 ) , .ZN( u2_u4_u0_n111 ) , .B1( u2_u4_u0_n118 ) , .A1( u2_u4_u0_n160 ) );
  INV_X1 u2_u4_u0_U3 (.A( u2_u4_u0_n113 ) , .ZN( u2_u4_u0_n166 ) );
  NAND2_X1 u2_u4_u0_U30 (.A1( u2_u4_u0_n100 ) , .ZN( u2_u4_u0_n129 ) , .A2( u2_u4_u0_n95 ) );
  INV_X1 u2_u4_u0_U31 (.A( u2_u4_u0_n118 ) , .ZN( u2_u4_u0_n158 ) );
  AOI21_X1 u2_u4_u0_U32 (.ZN( u2_u4_u0_n104 ) , .B1( u2_u4_u0_n107 ) , .B2( u2_u4_u0_n141 ) , .A( u2_u4_u0_n144 ) );
  AOI21_X1 u2_u4_u0_U33 (.B1( u2_u4_u0_n127 ) , .B2( u2_u4_u0_n129 ) , .A( u2_u4_u0_n138 ) , .ZN( u2_u4_u0_n96 ) );
  AOI21_X1 u2_u4_u0_U34 (.ZN( u2_u4_u0_n116 ) , .B2( u2_u4_u0_n142 ) , .A( u2_u4_u0_n144 ) , .B1( u2_u4_u0_n166 ) );
  NAND2_X1 u2_u4_u0_U35 (.A2( u2_u4_u0_n100 ) , .A1( u2_u4_u0_n101 ) , .ZN( u2_u4_u0_n139 ) );
  NAND2_X1 u2_u4_u0_U36 (.A2( u2_u4_u0_n100 ) , .ZN( u2_u4_u0_n131 ) , .A1( u2_u4_u0_n92 ) );
  NAND2_X1 u2_u4_u0_U37 (.A1( u2_u4_u0_n101 ) , .A2( u2_u4_u0_n102 ) , .ZN( u2_u4_u0_n150 ) );
  INV_X1 u2_u4_u0_U38 (.A( u2_u4_u0_n138 ) , .ZN( u2_u4_u0_n160 ) );
  NAND2_X1 u2_u4_u0_U39 (.A1( u2_u4_u0_n102 ) , .ZN( u2_u4_u0_n128 ) , .A2( u2_u4_u0_n95 ) );
  AOI21_X1 u2_u4_u0_U4 (.B1( u2_u4_u0_n114 ) , .ZN( u2_u4_u0_n115 ) , .B2( u2_u4_u0_n129 ) , .A( u2_u4_u0_n161 ) );
  NAND2_X1 u2_u4_u0_U40 (.ZN( u2_u4_u0_n148 ) , .A1( u2_u4_u0_n93 ) , .A2( u2_u4_u0_n95 ) );
  NAND2_X1 u2_u4_u0_U41 (.A2( u2_u4_u0_n102 ) , .A1( u2_u4_u0_n103 ) , .ZN( u2_u4_u0_n149 ) );
  NAND2_X1 u2_u4_u0_U42 (.A2( u2_u4_u0_n102 ) , .ZN( u2_u4_u0_n114 ) , .A1( u2_u4_u0_n92 ) );
  NAND2_X1 u2_u4_u0_U43 (.A2( u2_u4_u0_n101 ) , .ZN( u2_u4_u0_n121 ) , .A1( u2_u4_u0_n93 ) );
  NAND2_X1 u2_u4_u0_U44 (.ZN( u2_u4_u0_n112 ) , .A2( u2_u4_u0_n92 ) , .A1( u2_u4_u0_n93 ) );
  INV_X1 u2_u4_u0_U45 (.ZN( u2_u4_u0_n172 ) , .A( u2_u4_u0_n88 ) );
  OAI222_X1 u2_u4_u0_U46 (.C1( u2_u4_u0_n108 ) , .A1( u2_u4_u0_n125 ) , .B2( u2_u4_u0_n128 ) , .B1( u2_u4_u0_n144 ) , .A2( u2_u4_u0_n158 ) , .C2( u2_u4_u0_n161 ) , .ZN( u2_u4_u0_n88 ) );
  OR3_X1 u2_u4_u0_U47 (.A3( u2_u4_u0_n152 ) , .A2( u2_u4_u0_n153 ) , .A1( u2_u4_u0_n154 ) , .ZN( u2_u4_u0_n155 ) );
  AOI21_X1 u2_u4_u0_U48 (.B2( u2_u4_u0_n150 ) , .B1( u2_u4_u0_n151 ) , .ZN( u2_u4_u0_n152 ) , .A( u2_u4_u0_n158 ) );
  AOI21_X1 u2_u4_u0_U49 (.A( u2_u4_u0_n144 ) , .B2( u2_u4_u0_n145 ) , .B1( u2_u4_u0_n146 ) , .ZN( u2_u4_u0_n154 ) );
  AOI21_X1 u2_u4_u0_U5 (.B2( u2_u4_u0_n131 ) , .ZN( u2_u4_u0_n134 ) , .B1( u2_u4_u0_n151 ) , .A( u2_u4_u0_n158 ) );
  AOI21_X1 u2_u4_u0_U50 (.A( u2_u4_u0_n147 ) , .B2( u2_u4_u0_n148 ) , .B1( u2_u4_u0_n149 ) , .ZN( u2_u4_u0_n153 ) );
  INV_X1 u2_u4_u0_U51 (.ZN( u2_u4_u0_n171 ) , .A( u2_u4_u0_n99 ) );
  OAI211_X1 u2_u4_u0_U52 (.C2( u2_u4_u0_n140 ) , .C1( u2_u4_u0_n161 ) , .A( u2_u4_u0_n169 ) , .B( u2_u4_u0_n98 ) , .ZN( u2_u4_u0_n99 ) );
  AOI211_X1 u2_u4_u0_U53 (.C1( u2_u4_u0_n118 ) , .A( u2_u4_u0_n123 ) , .B( u2_u4_u0_n96 ) , .C2( u2_u4_u0_n97 ) , .ZN( u2_u4_u0_n98 ) );
  INV_X1 u2_u4_u0_U54 (.ZN( u2_u4_u0_n169 ) , .A( u2_u4_u0_n91 ) );
  NOR2_X1 u2_u4_u0_U55 (.A2( u2_u4_X_4 ) , .A1( u2_u4_X_5 ) , .ZN( u2_u4_u0_n118 ) );
  NOR2_X1 u2_u4_u0_U56 (.A2( u2_u4_X_2 ) , .ZN( u2_u4_u0_n103 ) , .A1( u2_u4_u0_n164 ) );
  NOR2_X1 u2_u4_u0_U57 (.A2( u2_u4_X_1 ) , .A1( u2_u4_X_2 ) , .ZN( u2_u4_u0_n92 ) );
  NOR2_X1 u2_u4_u0_U58 (.A2( u2_u4_X_1 ) , .ZN( u2_u4_u0_n101 ) , .A1( u2_u4_u0_n163 ) );
  NAND2_X1 u2_u4_u0_U59 (.A2( u2_u4_X_4 ) , .A1( u2_u4_X_5 ) , .ZN( u2_u4_u0_n144 ) );
  NOR2_X1 u2_u4_u0_U6 (.A1( u2_u4_u0_n108 ) , .ZN( u2_u4_u0_n123 ) , .A2( u2_u4_u0_n158 ) );
  NOR2_X1 u2_u4_u0_U60 (.A2( u2_u4_X_5 ) , .ZN( u2_u4_u0_n136 ) , .A1( u2_u4_u0_n159 ) );
  NAND2_X1 u2_u4_u0_U61 (.A1( u2_u4_X_5 ) , .ZN( u2_u4_u0_n138 ) , .A2( u2_u4_u0_n159 ) );
  AND2_X1 u2_u4_u0_U62 (.A2( u2_u4_X_3 ) , .A1( u2_u4_X_6 ) , .ZN( u2_u4_u0_n102 ) );
  INV_X1 u2_u4_u0_U63 (.A( u2_u4_X_4 ) , .ZN( u2_u4_u0_n159 ) );
  INV_X1 u2_u4_u0_U64 (.A( u2_u4_X_1 ) , .ZN( u2_u4_u0_n164 ) );
  INV_X1 u2_u4_u0_U65 (.A( u2_u4_X_2 ) , .ZN( u2_u4_u0_n163 ) );
  INV_X1 u2_u4_u0_U66 (.A( u2_u4_X_3 ) , .ZN( u2_u4_u0_n162 ) );
  AOI211_X1 u2_u4_u0_U67 (.B( u2_u4_u0_n133 ) , .A( u2_u4_u0_n134 ) , .C2( u2_u4_u0_n135 ) , .C1( u2_u4_u0_n136 ) , .ZN( u2_u4_u0_n137 ) );
  INV_X1 u2_u4_u0_U68 (.A( u2_u4_u0_n126 ) , .ZN( u2_u4_u0_n168 ) );
  INV_X1 u2_u4_u0_U69 (.ZN( u2_u4_u0_n174 ) , .A( u2_u4_u0_n89 ) );
  OAI21_X1 u2_u4_u0_U7 (.B1( u2_u4_u0_n150 ) , .B2( u2_u4_u0_n158 ) , .A( u2_u4_u0_n172 ) , .ZN( u2_u4_u0_n89 ) );
  AOI211_X1 u2_u4_u0_U70 (.B( u2_u4_u0_n104 ) , .A( u2_u4_u0_n105 ) , .ZN( u2_u4_u0_n106 ) , .C2( u2_u4_u0_n113 ) , .C1( u2_u4_u0_n160 ) );
  OR4_X1 u2_u4_u0_U71 (.ZN( u2_out4_31 ) , .A4( u2_u4_u0_n155 ) , .A2( u2_u4_u0_n156 ) , .A1( u2_u4_u0_n157 ) , .A3( u2_u4_u0_n173 ) );
  AOI21_X1 u2_u4_u0_U72 (.A( u2_u4_u0_n138 ) , .B2( u2_u4_u0_n139 ) , .B1( u2_u4_u0_n140 ) , .ZN( u2_u4_u0_n157 ) );
  AOI21_X1 u2_u4_u0_U73 (.B2( u2_u4_u0_n141 ) , .B1( u2_u4_u0_n142 ) , .ZN( u2_u4_u0_n156 ) , .A( u2_u4_u0_n161 ) );
  OR4_X1 u2_u4_u0_U74 (.ZN( u2_out4_17 ) , .A4( u2_u4_u0_n122 ) , .A2( u2_u4_u0_n123 ) , .A1( u2_u4_u0_n124 ) , .A3( u2_u4_u0_n170 ) );
  AOI21_X1 u2_u4_u0_U75 (.B2( u2_u4_u0_n107 ) , .ZN( u2_u4_u0_n124 ) , .B1( u2_u4_u0_n128 ) , .A( u2_u4_u0_n161 ) );
  INV_X1 u2_u4_u0_U76 (.A( u2_u4_u0_n111 ) , .ZN( u2_u4_u0_n170 ) );
  AOI21_X1 u2_u4_u0_U77 (.B1( u2_u4_u0_n132 ) , .ZN( u2_u4_u0_n133 ) , .A( u2_u4_u0_n144 ) , .B2( u2_u4_u0_n166 ) );
  OAI22_X1 u2_u4_u0_U78 (.ZN( u2_u4_u0_n105 ) , .A2( u2_u4_u0_n132 ) , .B1( u2_u4_u0_n146 ) , .A1( u2_u4_u0_n147 ) , .B2( u2_u4_u0_n161 ) );
  NAND2_X1 u2_u4_u0_U79 (.ZN( u2_u4_u0_n110 ) , .A2( u2_u4_u0_n132 ) , .A1( u2_u4_u0_n145 ) );
  AND2_X1 u2_u4_u0_U8 (.A1( u2_u4_u0_n114 ) , .A2( u2_u4_u0_n121 ) , .ZN( u2_u4_u0_n146 ) );
  INV_X1 u2_u4_u0_U80 (.A( u2_u4_u0_n119 ) , .ZN( u2_u4_u0_n167 ) );
  NAND2_X1 u2_u4_u0_U81 (.A2( u2_u4_u0_n103 ) , .ZN( u2_u4_u0_n140 ) , .A1( u2_u4_u0_n94 ) );
  NAND2_X1 u2_u4_u0_U82 (.A1( u2_u4_u0_n101 ) , .ZN( u2_u4_u0_n130 ) , .A2( u2_u4_u0_n94 ) );
  NAND2_X1 u2_u4_u0_U83 (.ZN( u2_u4_u0_n108 ) , .A1( u2_u4_u0_n92 ) , .A2( u2_u4_u0_n94 ) );
  AND2_X1 u2_u4_u0_U84 (.A1( u2_u4_X_6 ) , .A2( u2_u4_u0_n162 ) , .ZN( u2_u4_u0_n93 ) );
  NAND2_X1 u2_u4_u0_U85 (.ZN( u2_u4_u0_n142 ) , .A1( u2_u4_u0_n94 ) , .A2( u2_u4_u0_n95 ) );
  NOR2_X1 u2_u4_u0_U86 (.A2( u2_u4_X_6 ) , .ZN( u2_u4_u0_n100 ) , .A1( u2_u4_u0_n162 ) );
  NOR2_X1 u2_u4_u0_U87 (.A2( u2_u4_X_3 ) , .A1( u2_u4_X_6 ) , .ZN( u2_u4_u0_n94 ) );
  NAND3_X1 u2_u4_u0_U88 (.ZN( u2_out4_23 ) , .A3( u2_u4_u0_n137 ) , .A1( u2_u4_u0_n168 ) , .A2( u2_u4_u0_n171 ) );
  NAND3_X1 u2_u4_u0_U89 (.A3( u2_u4_u0_n127 ) , .A2( u2_u4_u0_n128 ) , .ZN( u2_u4_u0_n135 ) , .A1( u2_u4_u0_n150 ) );
  AND2_X1 u2_u4_u0_U9 (.A1( u2_u4_u0_n131 ) , .ZN( u2_u4_u0_n141 ) , .A2( u2_u4_u0_n150 ) );
  NAND3_X1 u2_u4_u0_U90 (.ZN( u2_u4_u0_n117 ) , .A3( u2_u4_u0_n132 ) , .A2( u2_u4_u0_n139 ) , .A1( u2_u4_u0_n148 ) );
  NAND3_X1 u2_u4_u0_U91 (.ZN( u2_u4_u0_n109 ) , .A2( u2_u4_u0_n114 ) , .A3( u2_u4_u0_n140 ) , .A1( u2_u4_u0_n149 ) );
  NAND3_X1 u2_u4_u0_U92 (.ZN( u2_out4_9 ) , .A3( u2_u4_u0_n106 ) , .A2( u2_u4_u0_n171 ) , .A1( u2_u4_u0_n174 ) );
  NAND3_X1 u2_u4_u0_U93 (.A2( u2_u4_u0_n128 ) , .A1( u2_u4_u0_n132 ) , .A3( u2_u4_u0_n146 ) , .ZN( u2_u4_u0_n97 ) );
  NOR2_X1 u2_u4_u1_U10 (.A1( u2_u4_u1_n112 ) , .A2( u2_u4_u1_n116 ) , .ZN( u2_u4_u1_n118 ) );
  NAND3_X1 u2_u4_u1_U100 (.ZN( u2_u4_u1_n113 ) , .A1( u2_u4_u1_n120 ) , .A3( u2_u4_u1_n133 ) , .A2( u2_u4_u1_n155 ) );
  OAI21_X1 u2_u4_u1_U11 (.ZN( u2_u4_u1_n101 ) , .B1( u2_u4_u1_n141 ) , .A( u2_u4_u1_n146 ) , .B2( u2_u4_u1_n183 ) );
  AOI21_X1 u2_u4_u1_U12 (.B2( u2_u4_u1_n155 ) , .B1( u2_u4_u1_n156 ) , .ZN( u2_u4_u1_n157 ) , .A( u2_u4_u1_n174 ) );
  NAND2_X1 u2_u4_u1_U13 (.ZN( u2_u4_u1_n140 ) , .A2( u2_u4_u1_n150 ) , .A1( u2_u4_u1_n155 ) );
  NAND2_X1 u2_u4_u1_U14 (.A1( u2_u4_u1_n131 ) , .ZN( u2_u4_u1_n147 ) , .A2( u2_u4_u1_n153 ) );
  INV_X1 u2_u4_u1_U15 (.A( u2_u4_u1_n139 ) , .ZN( u2_u4_u1_n174 ) );
  OR4_X1 u2_u4_u1_U16 (.A4( u2_u4_u1_n106 ) , .A3( u2_u4_u1_n107 ) , .ZN( u2_u4_u1_n108 ) , .A1( u2_u4_u1_n117 ) , .A2( u2_u4_u1_n184 ) );
  AOI21_X1 u2_u4_u1_U17 (.ZN( u2_u4_u1_n106 ) , .A( u2_u4_u1_n112 ) , .B1( u2_u4_u1_n154 ) , .B2( u2_u4_u1_n156 ) );
  AOI21_X1 u2_u4_u1_U18 (.ZN( u2_u4_u1_n107 ) , .B1( u2_u4_u1_n134 ) , .B2( u2_u4_u1_n149 ) , .A( u2_u4_u1_n174 ) );
  INV_X1 u2_u4_u1_U19 (.A( u2_u4_u1_n101 ) , .ZN( u2_u4_u1_n184 ) );
  INV_X1 u2_u4_u1_U20 (.A( u2_u4_u1_n112 ) , .ZN( u2_u4_u1_n171 ) );
  NAND2_X1 u2_u4_u1_U21 (.ZN( u2_u4_u1_n141 ) , .A1( u2_u4_u1_n153 ) , .A2( u2_u4_u1_n156 ) );
  AND2_X1 u2_u4_u1_U22 (.A1( u2_u4_u1_n123 ) , .ZN( u2_u4_u1_n134 ) , .A2( u2_u4_u1_n161 ) );
  NAND2_X1 u2_u4_u1_U23 (.A2( u2_u4_u1_n115 ) , .A1( u2_u4_u1_n116 ) , .ZN( u2_u4_u1_n148 ) );
  NAND2_X1 u2_u4_u1_U24 (.A2( u2_u4_u1_n133 ) , .A1( u2_u4_u1_n135 ) , .ZN( u2_u4_u1_n159 ) );
  NAND2_X1 u2_u4_u1_U25 (.A2( u2_u4_u1_n115 ) , .A1( u2_u4_u1_n120 ) , .ZN( u2_u4_u1_n132 ) );
  INV_X1 u2_u4_u1_U26 (.A( u2_u4_u1_n154 ) , .ZN( u2_u4_u1_n178 ) );
  INV_X1 u2_u4_u1_U27 (.A( u2_u4_u1_n151 ) , .ZN( u2_u4_u1_n183 ) );
  AND2_X1 u2_u4_u1_U28 (.A1( u2_u4_u1_n129 ) , .A2( u2_u4_u1_n133 ) , .ZN( u2_u4_u1_n149 ) );
  INV_X1 u2_u4_u1_U29 (.A( u2_u4_u1_n131 ) , .ZN( u2_u4_u1_n180 ) );
  INV_X1 u2_u4_u1_U3 (.A( u2_u4_u1_n159 ) , .ZN( u2_u4_u1_n182 ) );
  OAI221_X1 u2_u4_u1_U30 (.A( u2_u4_u1_n119 ) , .C2( u2_u4_u1_n129 ) , .ZN( u2_u4_u1_n138 ) , .B2( u2_u4_u1_n152 ) , .C1( u2_u4_u1_n174 ) , .B1( u2_u4_u1_n187 ) );
  INV_X1 u2_u4_u1_U31 (.A( u2_u4_u1_n148 ) , .ZN( u2_u4_u1_n187 ) );
  AOI211_X1 u2_u4_u1_U32 (.B( u2_u4_u1_n117 ) , .A( u2_u4_u1_n118 ) , .ZN( u2_u4_u1_n119 ) , .C2( u2_u4_u1_n146 ) , .C1( u2_u4_u1_n159 ) );
  NOR2_X1 u2_u4_u1_U33 (.A1( u2_u4_u1_n168 ) , .A2( u2_u4_u1_n176 ) , .ZN( u2_u4_u1_n98 ) );
  AOI211_X1 u2_u4_u1_U34 (.B( u2_u4_u1_n162 ) , .A( u2_u4_u1_n163 ) , .C2( u2_u4_u1_n164 ) , .ZN( u2_u4_u1_n165 ) , .C1( u2_u4_u1_n171 ) );
  AOI21_X1 u2_u4_u1_U35 (.A( u2_u4_u1_n160 ) , .B2( u2_u4_u1_n161 ) , .ZN( u2_u4_u1_n162 ) , .B1( u2_u4_u1_n182 ) );
  OR2_X1 u2_u4_u1_U36 (.A2( u2_u4_u1_n157 ) , .A1( u2_u4_u1_n158 ) , .ZN( u2_u4_u1_n163 ) );
  NAND2_X1 u2_u4_u1_U37 (.A1( u2_u4_u1_n128 ) , .ZN( u2_u4_u1_n146 ) , .A2( u2_u4_u1_n160 ) );
  NAND2_X1 u2_u4_u1_U38 (.A2( u2_u4_u1_n112 ) , .ZN( u2_u4_u1_n139 ) , .A1( u2_u4_u1_n152 ) );
  NAND2_X1 u2_u4_u1_U39 (.A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n156 ) , .A2( u2_u4_u1_n99 ) );
  AOI221_X1 u2_u4_u1_U4 (.A( u2_u4_u1_n138 ) , .C2( u2_u4_u1_n139 ) , .C1( u2_u4_u1_n140 ) , .B2( u2_u4_u1_n141 ) , .ZN( u2_u4_u1_n142 ) , .B1( u2_u4_u1_n175 ) );
  AOI221_X1 u2_u4_u1_U40 (.B1( u2_u4_u1_n140 ) , .ZN( u2_u4_u1_n167 ) , .B2( u2_u4_u1_n172 ) , .C2( u2_u4_u1_n175 ) , .C1( u2_u4_u1_n178 ) , .A( u2_u4_u1_n188 ) );
  INV_X1 u2_u4_u1_U41 (.ZN( u2_u4_u1_n188 ) , .A( u2_u4_u1_n97 ) );
  AOI211_X1 u2_u4_u1_U42 (.A( u2_u4_u1_n118 ) , .C1( u2_u4_u1_n132 ) , .C2( u2_u4_u1_n139 ) , .B( u2_u4_u1_n96 ) , .ZN( u2_u4_u1_n97 ) );
  AOI21_X1 u2_u4_u1_U43 (.B2( u2_u4_u1_n121 ) , .B1( u2_u4_u1_n135 ) , .A( u2_u4_u1_n152 ) , .ZN( u2_u4_u1_n96 ) );
  NOR2_X1 u2_u4_u1_U44 (.ZN( u2_u4_u1_n117 ) , .A1( u2_u4_u1_n121 ) , .A2( u2_u4_u1_n160 ) );
  OAI21_X1 u2_u4_u1_U45 (.B2( u2_u4_u1_n123 ) , .ZN( u2_u4_u1_n145 ) , .B1( u2_u4_u1_n160 ) , .A( u2_u4_u1_n185 ) );
  INV_X1 u2_u4_u1_U46 (.A( u2_u4_u1_n122 ) , .ZN( u2_u4_u1_n185 ) );
  AOI21_X1 u2_u4_u1_U47 (.B2( u2_u4_u1_n120 ) , .B1( u2_u4_u1_n121 ) , .ZN( u2_u4_u1_n122 ) , .A( u2_u4_u1_n128 ) );
  AOI21_X1 u2_u4_u1_U48 (.A( u2_u4_u1_n128 ) , .B2( u2_u4_u1_n129 ) , .ZN( u2_u4_u1_n130 ) , .B1( u2_u4_u1_n150 ) );
  NAND2_X1 u2_u4_u1_U49 (.ZN( u2_u4_u1_n112 ) , .A1( u2_u4_u1_n169 ) , .A2( u2_u4_u1_n170 ) );
  AOI211_X1 u2_u4_u1_U5 (.ZN( u2_u4_u1_n124 ) , .A( u2_u4_u1_n138 ) , .C2( u2_u4_u1_n139 ) , .B( u2_u4_u1_n145 ) , .C1( u2_u4_u1_n147 ) );
  NAND2_X1 u2_u4_u1_U50 (.ZN( u2_u4_u1_n129 ) , .A2( u2_u4_u1_n95 ) , .A1( u2_u4_u1_n98 ) );
  NAND2_X1 u2_u4_u1_U51 (.A1( u2_u4_u1_n102 ) , .ZN( u2_u4_u1_n154 ) , .A2( u2_u4_u1_n99 ) );
  NAND2_X1 u2_u4_u1_U52 (.A2( u2_u4_u1_n100 ) , .ZN( u2_u4_u1_n135 ) , .A1( u2_u4_u1_n99 ) );
  AOI21_X1 u2_u4_u1_U53 (.A( u2_u4_u1_n152 ) , .B2( u2_u4_u1_n153 ) , .B1( u2_u4_u1_n154 ) , .ZN( u2_u4_u1_n158 ) );
  INV_X1 u2_u4_u1_U54 (.A( u2_u4_u1_n160 ) , .ZN( u2_u4_u1_n175 ) );
  NAND2_X1 u2_u4_u1_U55 (.A1( u2_u4_u1_n100 ) , .ZN( u2_u4_u1_n116 ) , .A2( u2_u4_u1_n95 ) );
  NAND2_X1 u2_u4_u1_U56 (.A1( u2_u4_u1_n102 ) , .ZN( u2_u4_u1_n131 ) , .A2( u2_u4_u1_n95 ) );
  NAND2_X1 u2_u4_u1_U57 (.A2( u2_u4_u1_n104 ) , .ZN( u2_u4_u1_n121 ) , .A1( u2_u4_u1_n98 ) );
  NAND2_X1 u2_u4_u1_U58 (.A1( u2_u4_u1_n103 ) , .ZN( u2_u4_u1_n153 ) , .A2( u2_u4_u1_n98 ) );
  NAND2_X1 u2_u4_u1_U59 (.A2( u2_u4_u1_n104 ) , .A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n133 ) );
  AOI22_X1 u2_u4_u1_U6 (.B2( u2_u4_u1_n113 ) , .A2( u2_u4_u1_n114 ) , .ZN( u2_u4_u1_n125 ) , .A1( u2_u4_u1_n171 ) , .B1( u2_u4_u1_n173 ) );
  NAND2_X1 u2_u4_u1_U60 (.ZN( u2_u4_u1_n150 ) , .A2( u2_u4_u1_n98 ) , .A1( u2_u4_u1_n99 ) );
  NAND2_X1 u2_u4_u1_U61 (.A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n155 ) , .A2( u2_u4_u1_n95 ) );
  OAI21_X1 u2_u4_u1_U62 (.ZN( u2_u4_u1_n109 ) , .B1( u2_u4_u1_n129 ) , .B2( u2_u4_u1_n160 ) , .A( u2_u4_u1_n167 ) );
  NAND2_X1 u2_u4_u1_U63 (.A2( u2_u4_u1_n100 ) , .A1( u2_u4_u1_n103 ) , .ZN( u2_u4_u1_n120 ) );
  NAND2_X1 u2_u4_u1_U64 (.A1( u2_u4_u1_n102 ) , .A2( u2_u4_u1_n104 ) , .ZN( u2_u4_u1_n115 ) );
  NAND2_X1 u2_u4_u1_U65 (.A2( u2_u4_u1_n100 ) , .A1( u2_u4_u1_n104 ) , .ZN( u2_u4_u1_n151 ) );
  NAND2_X1 u2_u4_u1_U66 (.A2( u2_u4_u1_n103 ) , .A1( u2_u4_u1_n105 ) , .ZN( u2_u4_u1_n161 ) );
  INV_X1 u2_u4_u1_U67 (.A( u2_u4_u1_n152 ) , .ZN( u2_u4_u1_n173 ) );
  INV_X1 u2_u4_u1_U68 (.A( u2_u4_u1_n128 ) , .ZN( u2_u4_u1_n172 ) );
  NAND2_X1 u2_u4_u1_U69 (.A2( u2_u4_u1_n102 ) , .A1( u2_u4_u1_n103 ) , .ZN( u2_u4_u1_n123 ) );
  NAND2_X1 u2_u4_u1_U7 (.ZN( u2_u4_u1_n114 ) , .A1( u2_u4_u1_n134 ) , .A2( u2_u4_u1_n156 ) );
  NOR2_X1 u2_u4_u1_U70 (.A2( u2_u4_X_7 ) , .A1( u2_u4_X_8 ) , .ZN( u2_u4_u1_n95 ) );
  NOR2_X1 u2_u4_u1_U71 (.A1( u2_u4_X_12 ) , .A2( u2_u4_X_9 ) , .ZN( u2_u4_u1_n100 ) );
  NOR2_X1 u2_u4_u1_U72 (.A2( u2_u4_X_8 ) , .A1( u2_u4_u1_n177 ) , .ZN( u2_u4_u1_n99 ) );
  NOR2_X1 u2_u4_u1_U73 (.A2( u2_u4_X_12 ) , .ZN( u2_u4_u1_n102 ) , .A1( u2_u4_u1_n176 ) );
  NOR2_X1 u2_u4_u1_U74 (.A2( u2_u4_X_9 ) , .ZN( u2_u4_u1_n105 ) , .A1( u2_u4_u1_n168 ) );
  NAND2_X1 u2_u4_u1_U75 (.A1( u2_u4_X_10 ) , .ZN( u2_u4_u1_n160 ) , .A2( u2_u4_u1_n169 ) );
  NAND2_X1 u2_u4_u1_U76 (.A2( u2_u4_X_10 ) , .A1( u2_u4_X_11 ) , .ZN( u2_u4_u1_n152 ) );
  NAND2_X1 u2_u4_u1_U77 (.A1( u2_u4_X_11 ) , .ZN( u2_u4_u1_n128 ) , .A2( u2_u4_u1_n170 ) );
  AND2_X1 u2_u4_u1_U78 (.A2( u2_u4_X_7 ) , .A1( u2_u4_X_8 ) , .ZN( u2_u4_u1_n104 ) );
  AND2_X1 u2_u4_u1_U79 (.A1( u2_u4_X_8 ) , .ZN( u2_u4_u1_n103 ) , .A2( u2_u4_u1_n177 ) );
  AOI22_X1 u2_u4_u1_U8 (.B2( u2_u4_u1_n136 ) , .A2( u2_u4_u1_n137 ) , .ZN( u2_u4_u1_n143 ) , .A1( u2_u4_u1_n171 ) , .B1( u2_u4_u1_n173 ) );
  INV_X1 u2_u4_u1_U80 (.A( u2_u4_X_10 ) , .ZN( u2_u4_u1_n170 ) );
  INV_X1 u2_u4_u1_U81 (.A( u2_u4_X_9 ) , .ZN( u2_u4_u1_n176 ) );
  INV_X1 u2_u4_u1_U82 (.A( u2_u4_X_11 ) , .ZN( u2_u4_u1_n169 ) );
  INV_X1 u2_u4_u1_U83 (.A( u2_u4_X_12 ) , .ZN( u2_u4_u1_n168 ) );
  INV_X1 u2_u4_u1_U84 (.A( u2_u4_X_7 ) , .ZN( u2_u4_u1_n177 ) );
  NAND4_X1 u2_u4_u1_U85 (.ZN( u2_out4_28 ) , .A4( u2_u4_u1_n124 ) , .A3( u2_u4_u1_n125 ) , .A2( u2_u4_u1_n126 ) , .A1( u2_u4_u1_n127 ) );
  OAI21_X1 u2_u4_u1_U86 (.ZN( u2_u4_u1_n127 ) , .B2( u2_u4_u1_n139 ) , .B1( u2_u4_u1_n175 ) , .A( u2_u4_u1_n183 ) );
  OAI21_X1 u2_u4_u1_U87 (.ZN( u2_u4_u1_n126 ) , .B2( u2_u4_u1_n140 ) , .A( u2_u4_u1_n146 ) , .B1( u2_u4_u1_n178 ) );
  NAND4_X1 u2_u4_u1_U88 (.ZN( u2_out4_18 ) , .A4( u2_u4_u1_n165 ) , .A3( u2_u4_u1_n166 ) , .A1( u2_u4_u1_n167 ) , .A2( u2_u4_u1_n186 ) );
  AOI22_X1 u2_u4_u1_U89 (.B2( u2_u4_u1_n146 ) , .B1( u2_u4_u1_n147 ) , .A2( u2_u4_u1_n148 ) , .ZN( u2_u4_u1_n166 ) , .A1( u2_u4_u1_n172 ) );
  INV_X1 u2_u4_u1_U9 (.A( u2_u4_u1_n147 ) , .ZN( u2_u4_u1_n181 ) );
  INV_X1 u2_u4_u1_U90 (.A( u2_u4_u1_n145 ) , .ZN( u2_u4_u1_n186 ) );
  NAND4_X1 u2_u4_u1_U91 (.ZN( u2_out4_2 ) , .A4( u2_u4_u1_n142 ) , .A3( u2_u4_u1_n143 ) , .A2( u2_u4_u1_n144 ) , .A1( u2_u4_u1_n179 ) );
  OAI21_X1 u2_u4_u1_U92 (.B2( u2_u4_u1_n132 ) , .ZN( u2_u4_u1_n144 ) , .A( u2_u4_u1_n146 ) , .B1( u2_u4_u1_n180 ) );
  INV_X1 u2_u4_u1_U93 (.A( u2_u4_u1_n130 ) , .ZN( u2_u4_u1_n179 ) );
  OR4_X1 u2_u4_u1_U94 (.ZN( u2_out4_13 ) , .A4( u2_u4_u1_n108 ) , .A3( u2_u4_u1_n109 ) , .A2( u2_u4_u1_n110 ) , .A1( u2_u4_u1_n111 ) );
  AOI21_X1 u2_u4_u1_U95 (.ZN( u2_u4_u1_n111 ) , .A( u2_u4_u1_n128 ) , .B2( u2_u4_u1_n131 ) , .B1( u2_u4_u1_n135 ) );
  AOI21_X1 u2_u4_u1_U96 (.ZN( u2_u4_u1_n110 ) , .A( u2_u4_u1_n116 ) , .B1( u2_u4_u1_n152 ) , .B2( u2_u4_u1_n160 ) );
  NAND3_X1 u2_u4_u1_U97 (.A3( u2_u4_u1_n149 ) , .A2( u2_u4_u1_n150 ) , .A1( u2_u4_u1_n151 ) , .ZN( u2_u4_u1_n164 ) );
  NAND3_X1 u2_u4_u1_U98 (.A3( u2_u4_u1_n134 ) , .A2( u2_u4_u1_n135 ) , .ZN( u2_u4_u1_n136 ) , .A1( u2_u4_u1_n151 ) );
  NAND3_X1 u2_u4_u1_U99 (.A1( u2_u4_u1_n133 ) , .ZN( u2_u4_u1_n137 ) , .A2( u2_u4_u1_n154 ) , .A3( u2_u4_u1_n181 ) );
  OAI22_X1 u2_u4_u2_U10 (.ZN( u2_u4_u2_n109 ) , .A2( u2_u4_u2_n113 ) , .B2( u2_u4_u2_n133 ) , .B1( u2_u4_u2_n167 ) , .A1( u2_u4_u2_n168 ) );
  NAND3_X1 u2_u4_u2_U100 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n104 ) , .A3( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n98 ) );
  OAI22_X1 u2_u4_u2_U11 (.B1( u2_u4_u2_n151 ) , .A2( u2_u4_u2_n152 ) , .A1( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n160 ) , .B2( u2_u4_u2_n168 ) );
  NOR3_X1 u2_u4_u2_U12 (.A1( u2_u4_u2_n150 ) , .ZN( u2_u4_u2_n151 ) , .A3( u2_u4_u2_n175 ) , .A2( u2_u4_u2_n188 ) );
  AOI21_X1 u2_u4_u2_U13 (.ZN( u2_u4_u2_n144 ) , .B2( u2_u4_u2_n155 ) , .A( u2_u4_u2_n172 ) , .B1( u2_u4_u2_n185 ) );
  AOI21_X1 u2_u4_u2_U14 (.B2( u2_u4_u2_n143 ) , .ZN( u2_u4_u2_n145 ) , .B1( u2_u4_u2_n152 ) , .A( u2_u4_u2_n171 ) );
  AOI21_X1 u2_u4_u2_U15 (.B2( u2_u4_u2_n120 ) , .B1( u2_u4_u2_n121 ) , .ZN( u2_u4_u2_n126 ) , .A( u2_u4_u2_n167 ) );
  INV_X1 u2_u4_u2_U16 (.A( u2_u4_u2_n156 ) , .ZN( u2_u4_u2_n171 ) );
  INV_X1 u2_u4_u2_U17 (.A( u2_u4_u2_n120 ) , .ZN( u2_u4_u2_n188 ) );
  NAND2_X1 u2_u4_u2_U18 (.A2( u2_u4_u2_n122 ) , .ZN( u2_u4_u2_n150 ) , .A1( u2_u4_u2_n152 ) );
  INV_X1 u2_u4_u2_U19 (.A( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n170 ) );
  INV_X1 u2_u4_u2_U20 (.A( u2_u4_u2_n137 ) , .ZN( u2_u4_u2_n173 ) );
  NAND2_X1 u2_u4_u2_U21 (.A1( u2_u4_u2_n132 ) , .A2( u2_u4_u2_n139 ) , .ZN( u2_u4_u2_n157 ) );
  INV_X1 u2_u4_u2_U22 (.A( u2_u4_u2_n113 ) , .ZN( u2_u4_u2_n178 ) );
  INV_X1 u2_u4_u2_U23 (.A( u2_u4_u2_n139 ) , .ZN( u2_u4_u2_n175 ) );
  INV_X1 u2_u4_u2_U24 (.A( u2_u4_u2_n155 ) , .ZN( u2_u4_u2_n181 ) );
  INV_X1 u2_u4_u2_U25 (.A( u2_u4_u2_n119 ) , .ZN( u2_u4_u2_n177 ) );
  INV_X1 u2_u4_u2_U26 (.A( u2_u4_u2_n116 ) , .ZN( u2_u4_u2_n180 ) );
  INV_X1 u2_u4_u2_U27 (.A( u2_u4_u2_n131 ) , .ZN( u2_u4_u2_n179 ) );
  INV_X1 u2_u4_u2_U28 (.A( u2_u4_u2_n154 ) , .ZN( u2_u4_u2_n176 ) );
  NAND2_X1 u2_u4_u2_U29 (.A2( u2_u4_u2_n116 ) , .A1( u2_u4_u2_n117 ) , .ZN( u2_u4_u2_n118 ) );
  NOR2_X1 u2_u4_u2_U3 (.ZN( u2_u4_u2_n121 ) , .A2( u2_u4_u2_n177 ) , .A1( u2_u4_u2_n180 ) );
  INV_X1 u2_u4_u2_U30 (.A( u2_u4_u2_n132 ) , .ZN( u2_u4_u2_n182 ) );
  INV_X1 u2_u4_u2_U31 (.A( u2_u4_u2_n158 ) , .ZN( u2_u4_u2_n183 ) );
  OAI21_X1 u2_u4_u2_U32 (.A( u2_u4_u2_n156 ) , .B1( u2_u4_u2_n157 ) , .ZN( u2_u4_u2_n158 ) , .B2( u2_u4_u2_n179 ) );
  NOR2_X1 u2_u4_u2_U33 (.ZN( u2_u4_u2_n156 ) , .A1( u2_u4_u2_n166 ) , .A2( u2_u4_u2_n169 ) );
  NOR2_X1 u2_u4_u2_U34 (.A2( u2_u4_u2_n114 ) , .ZN( u2_u4_u2_n137 ) , .A1( u2_u4_u2_n140 ) );
  NOR2_X1 u2_u4_u2_U35 (.A2( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n153 ) , .A1( u2_u4_u2_n156 ) );
  AOI211_X1 u2_u4_u2_U36 (.ZN( u2_u4_u2_n130 ) , .C1( u2_u4_u2_n138 ) , .C2( u2_u4_u2_n179 ) , .B( u2_u4_u2_n96 ) , .A( u2_u4_u2_n97 ) );
  OAI22_X1 u2_u4_u2_U37 (.B1( u2_u4_u2_n133 ) , .A2( u2_u4_u2_n137 ) , .A1( u2_u4_u2_n152 ) , .B2( u2_u4_u2_n168 ) , .ZN( u2_u4_u2_n97 ) );
  OAI221_X1 u2_u4_u2_U38 (.B1( u2_u4_u2_n113 ) , .C1( u2_u4_u2_n132 ) , .A( u2_u4_u2_n149 ) , .B2( u2_u4_u2_n171 ) , .C2( u2_u4_u2_n172 ) , .ZN( u2_u4_u2_n96 ) );
  OAI221_X1 u2_u4_u2_U39 (.A( u2_u4_u2_n115 ) , .C2( u2_u4_u2_n123 ) , .B2( u2_u4_u2_n143 ) , .B1( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n163 ) , .C1( u2_u4_u2_n168 ) );
  INV_X1 u2_u4_u2_U4 (.A( u2_u4_u2_n134 ) , .ZN( u2_u4_u2_n185 ) );
  OAI21_X1 u2_u4_u2_U40 (.A( u2_u4_u2_n114 ) , .ZN( u2_u4_u2_n115 ) , .B1( u2_u4_u2_n176 ) , .B2( u2_u4_u2_n178 ) );
  OAI221_X1 u2_u4_u2_U41 (.A( u2_u4_u2_n135 ) , .B2( u2_u4_u2_n136 ) , .B1( u2_u4_u2_n137 ) , .ZN( u2_u4_u2_n162 ) , .C2( u2_u4_u2_n167 ) , .C1( u2_u4_u2_n185 ) );
  AND3_X1 u2_u4_u2_U42 (.A3( u2_u4_u2_n131 ) , .A2( u2_u4_u2_n132 ) , .A1( u2_u4_u2_n133 ) , .ZN( u2_u4_u2_n136 ) );
  AOI22_X1 u2_u4_u2_U43 (.ZN( u2_u4_u2_n135 ) , .B1( u2_u4_u2_n140 ) , .A1( u2_u4_u2_n156 ) , .B2( u2_u4_u2_n180 ) , .A2( u2_u4_u2_n188 ) );
  AOI21_X1 u2_u4_u2_U44 (.ZN( u2_u4_u2_n149 ) , .B1( u2_u4_u2_n173 ) , .B2( u2_u4_u2_n188 ) , .A( u2_u4_u2_n95 ) );
  AND3_X1 u2_u4_u2_U45 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n104 ) , .A3( u2_u4_u2_n156 ) , .ZN( u2_u4_u2_n95 ) );
  OAI21_X1 u2_u4_u2_U46 (.A( u2_u4_u2_n101 ) , .B2( u2_u4_u2_n121 ) , .B1( u2_u4_u2_n153 ) , .ZN( u2_u4_u2_n164 ) );
  NAND2_X1 u2_u4_u2_U47 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n107 ) , .ZN( u2_u4_u2_n155 ) );
  NAND2_X1 u2_u4_u2_U48 (.A2( u2_u4_u2_n105 ) , .A1( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n143 ) );
  NAND2_X1 u2_u4_u2_U49 (.A1( u2_u4_u2_n104 ) , .A2( u2_u4_u2_n106 ) , .ZN( u2_u4_u2_n152 ) );
  INV_X1 u2_u4_u2_U5 (.A( u2_u4_u2_n150 ) , .ZN( u2_u4_u2_n184 ) );
  NAND2_X1 u2_u4_u2_U50 (.A1( u2_u4_u2_n100 ) , .A2( u2_u4_u2_n105 ) , .ZN( u2_u4_u2_n132 ) );
  INV_X1 u2_u4_u2_U51 (.A( u2_u4_u2_n140 ) , .ZN( u2_u4_u2_n168 ) );
  INV_X1 u2_u4_u2_U52 (.A( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n167 ) );
  OAI21_X1 u2_u4_u2_U53 (.A( u2_u4_u2_n141 ) , .B2( u2_u4_u2_n142 ) , .ZN( u2_u4_u2_n146 ) , .B1( u2_u4_u2_n153 ) );
  OAI21_X1 u2_u4_u2_U54 (.A( u2_u4_u2_n140 ) , .ZN( u2_u4_u2_n141 ) , .B1( u2_u4_u2_n176 ) , .B2( u2_u4_u2_n177 ) );
  NOR3_X1 u2_u4_u2_U55 (.ZN( u2_u4_u2_n142 ) , .A3( u2_u4_u2_n175 ) , .A2( u2_u4_u2_n178 ) , .A1( u2_u4_u2_n181 ) );
  INV_X1 u2_u4_u2_U56 (.ZN( u2_u4_u2_n187 ) , .A( u2_u4_u2_n99 ) );
  OAI21_X1 u2_u4_u2_U57 (.B1( u2_u4_u2_n137 ) , .B2( u2_u4_u2_n143 ) , .A( u2_u4_u2_n98 ) , .ZN( u2_u4_u2_n99 ) );
  NAND2_X1 u2_u4_u2_U58 (.A1( u2_u4_u2_n102 ) , .A2( u2_u4_u2_n106 ) , .ZN( u2_u4_u2_n113 ) );
  NAND2_X1 u2_u4_u2_U59 (.A1( u2_u4_u2_n106 ) , .A2( u2_u4_u2_n107 ) , .ZN( u2_u4_u2_n131 ) );
  NOR4_X1 u2_u4_u2_U6 (.A4( u2_u4_u2_n124 ) , .A3( u2_u4_u2_n125 ) , .A2( u2_u4_u2_n126 ) , .A1( u2_u4_u2_n127 ) , .ZN( u2_u4_u2_n128 ) );
  NAND2_X1 u2_u4_u2_U60 (.A1( u2_u4_u2_n103 ) , .A2( u2_u4_u2_n107 ) , .ZN( u2_u4_u2_n139 ) );
  NAND2_X1 u2_u4_u2_U61 (.A1( u2_u4_u2_n103 ) , .A2( u2_u4_u2_n105 ) , .ZN( u2_u4_u2_n133 ) );
  NAND2_X1 u2_u4_u2_U62 (.A1( u2_u4_u2_n102 ) , .A2( u2_u4_u2_n103 ) , .ZN( u2_u4_u2_n154 ) );
  NAND2_X1 u2_u4_u2_U63 (.A2( u2_u4_u2_n103 ) , .A1( u2_u4_u2_n104 ) , .ZN( u2_u4_u2_n119 ) );
  NAND2_X1 u2_u4_u2_U64 (.A2( u2_u4_u2_n107 ) , .A1( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n123 ) );
  NAND2_X1 u2_u4_u2_U65 (.A1( u2_u4_u2_n104 ) , .A2( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n122 ) );
  INV_X1 u2_u4_u2_U66 (.A( u2_u4_u2_n114 ) , .ZN( u2_u4_u2_n172 ) );
  NAND2_X1 u2_u4_u2_U67 (.A2( u2_u4_u2_n100 ) , .A1( u2_u4_u2_n102 ) , .ZN( u2_u4_u2_n116 ) );
  NAND2_X1 u2_u4_u2_U68 (.A1( u2_u4_u2_n102 ) , .A2( u2_u4_u2_n108 ) , .ZN( u2_u4_u2_n120 ) );
  NAND2_X1 u2_u4_u2_U69 (.A2( u2_u4_u2_n105 ) , .A1( u2_u4_u2_n106 ) , .ZN( u2_u4_u2_n117 ) );
  AOI21_X1 u2_u4_u2_U7 (.B2( u2_u4_u2_n119 ) , .ZN( u2_u4_u2_n127 ) , .A( u2_u4_u2_n137 ) , .B1( u2_u4_u2_n155 ) );
  NOR2_X1 u2_u4_u2_U70 (.A2( u2_u4_X_16 ) , .ZN( u2_u4_u2_n140 ) , .A1( u2_u4_u2_n166 ) );
  NOR2_X1 u2_u4_u2_U71 (.A2( u2_u4_X_13 ) , .A1( u2_u4_X_14 ) , .ZN( u2_u4_u2_n100 ) );
  NOR2_X1 u2_u4_u2_U72 (.A2( u2_u4_X_16 ) , .A1( u2_u4_X_17 ) , .ZN( u2_u4_u2_n138 ) );
  NOR2_X1 u2_u4_u2_U73 (.A2( u2_u4_X_15 ) , .A1( u2_u4_X_18 ) , .ZN( u2_u4_u2_n104 ) );
  NOR2_X1 u2_u4_u2_U74 (.A2( u2_u4_X_14 ) , .ZN( u2_u4_u2_n103 ) , .A1( u2_u4_u2_n174 ) );
  NOR2_X1 u2_u4_u2_U75 (.A2( u2_u4_X_15 ) , .ZN( u2_u4_u2_n102 ) , .A1( u2_u4_u2_n165 ) );
  NOR2_X1 u2_u4_u2_U76 (.A2( u2_u4_X_17 ) , .ZN( u2_u4_u2_n114 ) , .A1( u2_u4_u2_n169 ) );
  AND2_X1 u2_u4_u2_U77 (.A1( u2_u4_X_15 ) , .ZN( u2_u4_u2_n105 ) , .A2( u2_u4_u2_n165 ) );
  AND2_X1 u2_u4_u2_U78 (.A2( u2_u4_X_15 ) , .A1( u2_u4_X_18 ) , .ZN( u2_u4_u2_n107 ) );
  AND2_X1 u2_u4_u2_U79 (.A1( u2_u4_X_14 ) , .ZN( u2_u4_u2_n106 ) , .A2( u2_u4_u2_n174 ) );
  AOI21_X1 u2_u4_u2_U8 (.ZN( u2_u4_u2_n124 ) , .B1( u2_u4_u2_n131 ) , .B2( u2_u4_u2_n143 ) , .A( u2_u4_u2_n172 ) );
  AND2_X1 u2_u4_u2_U80 (.A1( u2_u4_X_13 ) , .A2( u2_u4_X_14 ) , .ZN( u2_u4_u2_n108 ) );
  INV_X1 u2_u4_u2_U81 (.A( u2_u4_X_16 ) , .ZN( u2_u4_u2_n169 ) );
  INV_X1 u2_u4_u2_U82 (.A( u2_u4_X_17 ) , .ZN( u2_u4_u2_n166 ) );
  INV_X1 u2_u4_u2_U83 (.A( u2_u4_X_13 ) , .ZN( u2_u4_u2_n174 ) );
  INV_X1 u2_u4_u2_U84 (.A( u2_u4_X_18 ) , .ZN( u2_u4_u2_n165 ) );
  NAND4_X1 u2_u4_u2_U85 (.ZN( u2_out4_30 ) , .A4( u2_u4_u2_n147 ) , .A3( u2_u4_u2_n148 ) , .A2( u2_u4_u2_n149 ) , .A1( u2_u4_u2_n187 ) );
  NOR3_X1 u2_u4_u2_U86 (.A3( u2_u4_u2_n144 ) , .A2( u2_u4_u2_n145 ) , .A1( u2_u4_u2_n146 ) , .ZN( u2_u4_u2_n147 ) );
  AOI21_X1 u2_u4_u2_U87 (.B2( u2_u4_u2_n138 ) , .ZN( u2_u4_u2_n148 ) , .A( u2_u4_u2_n162 ) , .B1( u2_u4_u2_n182 ) );
  NAND4_X1 u2_u4_u2_U88 (.ZN( u2_out4_24 ) , .A4( u2_u4_u2_n111 ) , .A3( u2_u4_u2_n112 ) , .A1( u2_u4_u2_n130 ) , .A2( u2_u4_u2_n187 ) );
  AOI221_X1 u2_u4_u2_U89 (.A( u2_u4_u2_n109 ) , .B1( u2_u4_u2_n110 ) , .ZN( u2_u4_u2_n111 ) , .C1( u2_u4_u2_n134 ) , .C2( u2_u4_u2_n170 ) , .B2( u2_u4_u2_n173 ) );
  AOI21_X1 u2_u4_u2_U9 (.B2( u2_u4_u2_n123 ) , .ZN( u2_u4_u2_n125 ) , .A( u2_u4_u2_n171 ) , .B1( u2_u4_u2_n184 ) );
  AOI21_X1 u2_u4_u2_U90 (.ZN( u2_u4_u2_n112 ) , .B2( u2_u4_u2_n156 ) , .A( u2_u4_u2_n164 ) , .B1( u2_u4_u2_n181 ) );
  NAND4_X1 u2_u4_u2_U91 (.ZN( u2_out4_16 ) , .A4( u2_u4_u2_n128 ) , .A3( u2_u4_u2_n129 ) , .A1( u2_u4_u2_n130 ) , .A2( u2_u4_u2_n186 ) );
  AOI22_X1 u2_u4_u2_U92 (.A2( u2_u4_u2_n118 ) , .ZN( u2_u4_u2_n129 ) , .A1( u2_u4_u2_n140 ) , .B1( u2_u4_u2_n157 ) , .B2( u2_u4_u2_n170 ) );
  INV_X1 u2_u4_u2_U93 (.A( u2_u4_u2_n163 ) , .ZN( u2_u4_u2_n186 ) );
  OR4_X1 u2_u4_u2_U94 (.ZN( u2_out4_6 ) , .A4( u2_u4_u2_n161 ) , .A3( u2_u4_u2_n162 ) , .A2( u2_u4_u2_n163 ) , .A1( u2_u4_u2_n164 ) );
  OR3_X1 u2_u4_u2_U95 (.A2( u2_u4_u2_n159 ) , .A1( u2_u4_u2_n160 ) , .ZN( u2_u4_u2_n161 ) , .A3( u2_u4_u2_n183 ) );
  AOI21_X1 u2_u4_u2_U96 (.B2( u2_u4_u2_n154 ) , .B1( u2_u4_u2_n155 ) , .ZN( u2_u4_u2_n159 ) , .A( u2_u4_u2_n167 ) );
  NAND3_X1 u2_u4_u2_U97 (.A2( u2_u4_u2_n117 ) , .A1( u2_u4_u2_n122 ) , .A3( u2_u4_u2_n123 ) , .ZN( u2_u4_u2_n134 ) );
  NAND3_X1 u2_u4_u2_U98 (.ZN( u2_u4_u2_n110 ) , .A2( u2_u4_u2_n131 ) , .A3( u2_u4_u2_n139 ) , .A1( u2_u4_u2_n154 ) );
  NAND3_X1 u2_u4_u2_U99 (.A2( u2_u4_u2_n100 ) , .ZN( u2_u4_u2_n101 ) , .A1( u2_u4_u2_n104 ) , .A3( u2_u4_u2_n114 ) );
  OAI22_X1 u2_u4_u3_U10 (.B1( u2_u4_u3_n113 ) , .A2( u2_u4_u3_n135 ) , .A1( u2_u4_u3_n150 ) , .B2( u2_u4_u3_n164 ) , .ZN( u2_u4_u3_n98 ) );
  OAI211_X1 u2_u4_u3_U11 (.B( u2_u4_u3_n106 ) , .ZN( u2_u4_u3_n119 ) , .C2( u2_u4_u3_n128 ) , .C1( u2_u4_u3_n167 ) , .A( u2_u4_u3_n181 ) );
  AOI221_X1 u2_u4_u3_U12 (.C1( u2_u4_u3_n105 ) , .ZN( u2_u4_u3_n106 ) , .A( u2_u4_u3_n131 ) , .B2( u2_u4_u3_n132 ) , .C2( u2_u4_u3_n133 ) , .B1( u2_u4_u3_n169 ) );
  INV_X1 u2_u4_u3_U13 (.ZN( u2_u4_u3_n181 ) , .A( u2_u4_u3_n98 ) );
  NAND2_X1 u2_u4_u3_U14 (.ZN( u2_u4_u3_n105 ) , .A2( u2_u4_u3_n130 ) , .A1( u2_u4_u3_n155 ) );
  AOI22_X1 u2_u4_u3_U15 (.B1( u2_u4_u3_n115 ) , .A2( u2_u4_u3_n116 ) , .ZN( u2_u4_u3_n123 ) , .B2( u2_u4_u3_n133 ) , .A1( u2_u4_u3_n169 ) );
  NAND2_X1 u2_u4_u3_U16 (.ZN( u2_u4_u3_n116 ) , .A2( u2_u4_u3_n151 ) , .A1( u2_u4_u3_n182 ) );
  NOR2_X1 u2_u4_u3_U17 (.ZN( u2_u4_u3_n126 ) , .A2( u2_u4_u3_n150 ) , .A1( u2_u4_u3_n164 ) );
  AOI21_X1 u2_u4_u3_U18 (.ZN( u2_u4_u3_n112 ) , .B2( u2_u4_u3_n146 ) , .B1( u2_u4_u3_n155 ) , .A( u2_u4_u3_n167 ) );
  NAND2_X1 u2_u4_u3_U19 (.A1( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n142 ) , .A2( u2_u4_u3_n164 ) );
  NAND2_X1 u2_u4_u3_U20 (.ZN( u2_u4_u3_n132 ) , .A2( u2_u4_u3_n152 ) , .A1( u2_u4_u3_n156 ) );
  AND2_X1 u2_u4_u3_U21 (.A2( u2_u4_u3_n113 ) , .A1( u2_u4_u3_n114 ) , .ZN( u2_u4_u3_n151 ) );
  INV_X1 u2_u4_u3_U22 (.A( u2_u4_u3_n133 ) , .ZN( u2_u4_u3_n165 ) );
  INV_X1 u2_u4_u3_U23 (.A( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n170 ) );
  NAND2_X1 u2_u4_u3_U24 (.A1( u2_u4_u3_n107 ) , .A2( u2_u4_u3_n108 ) , .ZN( u2_u4_u3_n140 ) );
  NAND2_X1 u2_u4_u3_U25 (.ZN( u2_u4_u3_n117 ) , .A1( u2_u4_u3_n124 ) , .A2( u2_u4_u3_n148 ) );
  NAND2_X1 u2_u4_u3_U26 (.ZN( u2_u4_u3_n143 ) , .A1( u2_u4_u3_n165 ) , .A2( u2_u4_u3_n167 ) );
  INV_X1 u2_u4_u3_U27 (.A( u2_u4_u3_n130 ) , .ZN( u2_u4_u3_n177 ) );
  INV_X1 u2_u4_u3_U28 (.A( u2_u4_u3_n128 ) , .ZN( u2_u4_u3_n176 ) );
  INV_X1 u2_u4_u3_U29 (.A( u2_u4_u3_n155 ) , .ZN( u2_u4_u3_n174 ) );
  INV_X1 u2_u4_u3_U3 (.A( u2_u4_u3_n129 ) , .ZN( u2_u4_u3_n183 ) );
  INV_X1 u2_u4_u3_U30 (.A( u2_u4_u3_n139 ) , .ZN( u2_u4_u3_n185 ) );
  NOR2_X1 u2_u4_u3_U31 (.ZN( u2_u4_u3_n135 ) , .A2( u2_u4_u3_n141 ) , .A1( u2_u4_u3_n169 ) );
  OAI222_X1 u2_u4_u3_U32 (.C2( u2_u4_u3_n107 ) , .A2( u2_u4_u3_n108 ) , .B1( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n138 ) , .B2( u2_u4_u3_n146 ) , .C1( u2_u4_u3_n154 ) , .A1( u2_u4_u3_n164 ) );
  NOR4_X1 u2_u4_u3_U33 (.A4( u2_u4_u3_n157 ) , .A3( u2_u4_u3_n158 ) , .A2( u2_u4_u3_n159 ) , .A1( u2_u4_u3_n160 ) , .ZN( u2_u4_u3_n161 ) );
  AOI21_X1 u2_u4_u3_U34 (.B2( u2_u4_u3_n152 ) , .B1( u2_u4_u3_n153 ) , .ZN( u2_u4_u3_n158 ) , .A( u2_u4_u3_n164 ) );
  AOI21_X1 u2_u4_u3_U35 (.A( u2_u4_u3_n149 ) , .B2( u2_u4_u3_n150 ) , .B1( u2_u4_u3_n151 ) , .ZN( u2_u4_u3_n159 ) );
  AOI21_X1 u2_u4_u3_U36 (.A( u2_u4_u3_n154 ) , .B2( u2_u4_u3_n155 ) , .B1( u2_u4_u3_n156 ) , .ZN( u2_u4_u3_n157 ) );
  AOI211_X1 u2_u4_u3_U37 (.ZN( u2_u4_u3_n109 ) , .A( u2_u4_u3_n119 ) , .C2( u2_u4_u3_n129 ) , .B( u2_u4_u3_n138 ) , .C1( u2_u4_u3_n141 ) );
  AOI211_X1 u2_u4_u3_U38 (.B( u2_u4_u3_n119 ) , .A( u2_u4_u3_n120 ) , .C2( u2_u4_u3_n121 ) , .ZN( u2_u4_u3_n122 ) , .C1( u2_u4_u3_n179 ) );
  INV_X1 u2_u4_u3_U39 (.A( u2_u4_u3_n156 ) , .ZN( u2_u4_u3_n179 ) );
  INV_X1 u2_u4_u3_U4 (.A( u2_u4_u3_n140 ) , .ZN( u2_u4_u3_n182 ) );
  OAI22_X1 u2_u4_u3_U40 (.B1( u2_u4_u3_n118 ) , .ZN( u2_u4_u3_n120 ) , .A1( u2_u4_u3_n135 ) , .B2( u2_u4_u3_n154 ) , .A2( u2_u4_u3_n178 ) );
  AND3_X1 u2_u4_u3_U41 (.ZN( u2_u4_u3_n118 ) , .A2( u2_u4_u3_n124 ) , .A1( u2_u4_u3_n144 ) , .A3( u2_u4_u3_n152 ) );
  INV_X1 u2_u4_u3_U42 (.A( u2_u4_u3_n121 ) , .ZN( u2_u4_u3_n164 ) );
  NAND2_X1 u2_u4_u3_U43 (.ZN( u2_u4_u3_n133 ) , .A1( u2_u4_u3_n154 ) , .A2( u2_u4_u3_n164 ) );
  OAI211_X1 u2_u4_u3_U44 (.B( u2_u4_u3_n127 ) , .ZN( u2_u4_u3_n139 ) , .C1( u2_u4_u3_n150 ) , .C2( u2_u4_u3_n154 ) , .A( u2_u4_u3_n184 ) );
  INV_X1 u2_u4_u3_U45 (.A( u2_u4_u3_n125 ) , .ZN( u2_u4_u3_n184 ) );
  AOI221_X1 u2_u4_u3_U46 (.A( u2_u4_u3_n126 ) , .ZN( u2_u4_u3_n127 ) , .C2( u2_u4_u3_n132 ) , .C1( u2_u4_u3_n169 ) , .B2( u2_u4_u3_n170 ) , .B1( u2_u4_u3_n174 ) );
  OAI22_X1 u2_u4_u3_U47 (.A1( u2_u4_u3_n124 ) , .ZN( u2_u4_u3_n125 ) , .B2( u2_u4_u3_n145 ) , .A2( u2_u4_u3_n165 ) , .B1( u2_u4_u3_n167 ) );
  NOR2_X1 u2_u4_u3_U48 (.A1( u2_u4_u3_n113 ) , .ZN( u2_u4_u3_n131 ) , .A2( u2_u4_u3_n154 ) );
  NAND2_X1 u2_u4_u3_U49 (.A1( u2_u4_u3_n103 ) , .ZN( u2_u4_u3_n150 ) , .A2( u2_u4_u3_n99 ) );
  INV_X1 u2_u4_u3_U5 (.A( u2_u4_u3_n117 ) , .ZN( u2_u4_u3_n178 ) );
  NAND2_X1 u2_u4_u3_U50 (.A2( u2_u4_u3_n102 ) , .ZN( u2_u4_u3_n155 ) , .A1( u2_u4_u3_n97 ) );
  INV_X1 u2_u4_u3_U51 (.A( u2_u4_u3_n141 ) , .ZN( u2_u4_u3_n167 ) );
  AOI21_X1 u2_u4_u3_U52 (.B2( u2_u4_u3_n114 ) , .B1( u2_u4_u3_n146 ) , .A( u2_u4_u3_n154 ) , .ZN( u2_u4_u3_n94 ) );
  AOI21_X1 u2_u4_u3_U53 (.ZN( u2_u4_u3_n110 ) , .B2( u2_u4_u3_n142 ) , .B1( u2_u4_u3_n186 ) , .A( u2_u4_u3_n95 ) );
  INV_X1 u2_u4_u3_U54 (.A( u2_u4_u3_n145 ) , .ZN( u2_u4_u3_n186 ) );
  AOI21_X1 u2_u4_u3_U55 (.B1( u2_u4_u3_n124 ) , .A( u2_u4_u3_n149 ) , .B2( u2_u4_u3_n155 ) , .ZN( u2_u4_u3_n95 ) );
  INV_X1 u2_u4_u3_U56 (.A( u2_u4_u3_n149 ) , .ZN( u2_u4_u3_n169 ) );
  NAND2_X1 u2_u4_u3_U57 (.ZN( u2_u4_u3_n124 ) , .A1( u2_u4_u3_n96 ) , .A2( u2_u4_u3_n97 ) );
  NAND2_X1 u2_u4_u3_U58 (.A2( u2_u4_u3_n100 ) , .ZN( u2_u4_u3_n146 ) , .A1( u2_u4_u3_n96 ) );
  NAND2_X1 u2_u4_u3_U59 (.A1( u2_u4_u3_n101 ) , .ZN( u2_u4_u3_n145 ) , .A2( u2_u4_u3_n99 ) );
  AOI221_X1 u2_u4_u3_U6 (.A( u2_u4_u3_n131 ) , .C2( u2_u4_u3_n132 ) , .C1( u2_u4_u3_n133 ) , .ZN( u2_u4_u3_n134 ) , .B1( u2_u4_u3_n143 ) , .B2( u2_u4_u3_n177 ) );
  NAND2_X1 u2_u4_u3_U60 (.A1( u2_u4_u3_n100 ) , .ZN( u2_u4_u3_n156 ) , .A2( u2_u4_u3_n99 ) );
  NAND2_X1 u2_u4_u3_U61 (.A2( u2_u4_u3_n101 ) , .A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n148 ) );
  NAND2_X1 u2_u4_u3_U62 (.A1( u2_u4_u3_n100 ) , .A2( u2_u4_u3_n102 ) , .ZN( u2_u4_u3_n128 ) );
  NAND2_X1 u2_u4_u3_U63 (.A2( u2_u4_u3_n101 ) , .A1( u2_u4_u3_n102 ) , .ZN( u2_u4_u3_n152 ) );
  NAND2_X1 u2_u4_u3_U64 (.A2( u2_u4_u3_n101 ) , .ZN( u2_u4_u3_n114 ) , .A1( u2_u4_u3_n96 ) );
  NAND2_X1 u2_u4_u3_U65 (.ZN( u2_u4_u3_n107 ) , .A1( u2_u4_u3_n97 ) , .A2( u2_u4_u3_n99 ) );
  NAND2_X1 u2_u4_u3_U66 (.A2( u2_u4_u3_n100 ) , .A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n113 ) );
  NAND2_X1 u2_u4_u3_U67 (.A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n153 ) , .A2( u2_u4_u3_n97 ) );
  NAND2_X1 u2_u4_u3_U68 (.A2( u2_u4_u3_n103 ) , .A1( u2_u4_u3_n104 ) , .ZN( u2_u4_u3_n130 ) );
  NAND2_X1 u2_u4_u3_U69 (.A2( u2_u4_u3_n103 ) , .ZN( u2_u4_u3_n144 ) , .A1( u2_u4_u3_n96 ) );
  OAI22_X1 u2_u4_u3_U7 (.B2( u2_u4_u3_n147 ) , .A2( u2_u4_u3_n148 ) , .ZN( u2_u4_u3_n160 ) , .B1( u2_u4_u3_n165 ) , .A1( u2_u4_u3_n168 ) );
  NAND2_X1 u2_u4_u3_U70 (.A1( u2_u4_u3_n102 ) , .A2( u2_u4_u3_n103 ) , .ZN( u2_u4_u3_n108 ) );
  NOR2_X1 u2_u4_u3_U71 (.A2( u2_u4_X_19 ) , .A1( u2_u4_X_20 ) , .ZN( u2_u4_u3_n99 ) );
  NOR2_X1 u2_u4_u3_U72 (.A2( u2_u4_X_21 ) , .A1( u2_u4_X_24 ) , .ZN( u2_u4_u3_n103 ) );
  NOR2_X1 u2_u4_u3_U73 (.A2( u2_u4_X_24 ) , .A1( u2_u4_u3_n171 ) , .ZN( u2_u4_u3_n97 ) );
  NOR2_X1 u2_u4_u3_U74 (.A2( u2_u4_X_23 ) , .ZN( u2_u4_u3_n141 ) , .A1( u2_u4_u3_n166 ) );
  NOR2_X1 u2_u4_u3_U75 (.A2( u2_u4_X_19 ) , .A1( u2_u4_u3_n172 ) , .ZN( u2_u4_u3_n96 ) );
  NAND2_X1 u2_u4_u3_U76 (.A1( u2_u4_X_22 ) , .A2( u2_u4_X_23 ) , .ZN( u2_u4_u3_n154 ) );
  NAND2_X1 u2_u4_u3_U77 (.A1( u2_u4_X_23 ) , .ZN( u2_u4_u3_n149 ) , .A2( u2_u4_u3_n166 ) );
  NOR2_X1 u2_u4_u3_U78 (.A2( u2_u4_X_22 ) , .A1( u2_u4_X_23 ) , .ZN( u2_u4_u3_n121 ) );
  AND2_X1 u2_u4_u3_U79 (.A1( u2_u4_X_24 ) , .ZN( u2_u4_u3_n101 ) , .A2( u2_u4_u3_n171 ) );
  AND3_X1 u2_u4_u3_U8 (.A3( u2_u4_u3_n144 ) , .A2( u2_u4_u3_n145 ) , .A1( u2_u4_u3_n146 ) , .ZN( u2_u4_u3_n147 ) );
  AND2_X1 u2_u4_u3_U80 (.A1( u2_u4_X_19 ) , .ZN( u2_u4_u3_n102 ) , .A2( u2_u4_u3_n172 ) );
  AND2_X1 u2_u4_u3_U81 (.A1( u2_u4_X_21 ) , .A2( u2_u4_X_24 ) , .ZN( u2_u4_u3_n100 ) );
  AND2_X1 u2_u4_u3_U82 (.A2( u2_u4_X_19 ) , .A1( u2_u4_X_20 ) , .ZN( u2_u4_u3_n104 ) );
  INV_X1 u2_u4_u3_U83 (.A( u2_u4_X_22 ) , .ZN( u2_u4_u3_n166 ) );
  INV_X1 u2_u4_u3_U84 (.A( u2_u4_X_21 ) , .ZN( u2_u4_u3_n171 ) );
  INV_X1 u2_u4_u3_U85 (.A( u2_u4_X_20 ) , .ZN( u2_u4_u3_n172 ) );
  OR4_X1 u2_u4_u3_U86 (.ZN( u2_out4_10 ) , .A4( u2_u4_u3_n136 ) , .A3( u2_u4_u3_n137 ) , .A1( u2_u4_u3_n138 ) , .A2( u2_u4_u3_n139 ) );
  OAI222_X1 u2_u4_u3_U87 (.C1( u2_u4_u3_n128 ) , .ZN( u2_u4_u3_n137 ) , .B1( u2_u4_u3_n148 ) , .A2( u2_u4_u3_n150 ) , .B2( u2_u4_u3_n154 ) , .C2( u2_u4_u3_n164 ) , .A1( u2_u4_u3_n167 ) );
  OAI221_X1 u2_u4_u3_U88 (.A( u2_u4_u3_n134 ) , .B2( u2_u4_u3_n135 ) , .ZN( u2_u4_u3_n136 ) , .C1( u2_u4_u3_n149 ) , .B1( u2_u4_u3_n151 ) , .C2( u2_u4_u3_n183 ) );
  NAND4_X1 u2_u4_u3_U89 (.ZN( u2_out4_26 ) , .A4( u2_u4_u3_n109 ) , .A3( u2_u4_u3_n110 ) , .A2( u2_u4_u3_n111 ) , .A1( u2_u4_u3_n173 ) );
  INV_X1 u2_u4_u3_U9 (.A( u2_u4_u3_n143 ) , .ZN( u2_u4_u3_n168 ) );
  INV_X1 u2_u4_u3_U90 (.ZN( u2_u4_u3_n173 ) , .A( u2_u4_u3_n94 ) );
  OAI21_X1 u2_u4_u3_U91 (.ZN( u2_u4_u3_n111 ) , .B2( u2_u4_u3_n117 ) , .A( u2_u4_u3_n133 ) , .B1( u2_u4_u3_n176 ) );
  NAND4_X1 u2_u4_u3_U92 (.ZN( u2_out4_20 ) , .A4( u2_u4_u3_n122 ) , .A3( u2_u4_u3_n123 ) , .A1( u2_u4_u3_n175 ) , .A2( u2_u4_u3_n180 ) );
  INV_X1 u2_u4_u3_U93 (.A( u2_u4_u3_n126 ) , .ZN( u2_u4_u3_n180 ) );
  INV_X1 u2_u4_u3_U94 (.A( u2_u4_u3_n112 ) , .ZN( u2_u4_u3_n175 ) );
  NAND4_X1 u2_u4_u3_U95 (.ZN( u2_out4_1 ) , .A4( u2_u4_u3_n161 ) , .A3( u2_u4_u3_n162 ) , .A2( u2_u4_u3_n163 ) , .A1( u2_u4_u3_n185 ) );
  NAND2_X1 u2_u4_u3_U96 (.ZN( u2_u4_u3_n163 ) , .A2( u2_u4_u3_n170 ) , .A1( u2_u4_u3_n176 ) );
  AOI22_X1 u2_u4_u3_U97 (.B2( u2_u4_u3_n140 ) , .B1( u2_u4_u3_n141 ) , .A2( u2_u4_u3_n142 ) , .ZN( u2_u4_u3_n162 ) , .A1( u2_u4_u3_n177 ) );
  NAND3_X1 u2_u4_u3_U98 (.A1( u2_u4_u3_n114 ) , .ZN( u2_u4_u3_n115 ) , .A2( u2_u4_u3_n145 ) , .A3( u2_u4_u3_n153 ) );
  NAND3_X1 u2_u4_u3_U99 (.ZN( u2_u4_u3_n129 ) , .A2( u2_u4_u3_n144 ) , .A1( u2_u4_u3_n153 ) , .A3( u2_u4_u3_n182 ) );
  OAI22_X1 u2_u4_u4_U10 (.B2( u2_u4_u4_n135 ) , .ZN( u2_u4_u4_n137 ) , .B1( u2_u4_u4_n153 ) , .A1( u2_u4_u4_n155 ) , .A2( u2_u4_u4_n171 ) );
  AND3_X1 u2_u4_u4_U11 (.A2( u2_u4_u4_n134 ) , .ZN( u2_u4_u4_n135 ) , .A3( u2_u4_u4_n145 ) , .A1( u2_u4_u4_n157 ) );
  NAND2_X1 u2_u4_u4_U12 (.ZN( u2_u4_u4_n132 ) , .A2( u2_u4_u4_n170 ) , .A1( u2_u4_u4_n173 ) );
  AOI21_X1 u2_u4_u4_U13 (.B2( u2_u4_u4_n160 ) , .B1( u2_u4_u4_n161 ) , .ZN( u2_u4_u4_n162 ) , .A( u2_u4_u4_n170 ) );
  AOI21_X1 u2_u4_u4_U14 (.ZN( u2_u4_u4_n107 ) , .B2( u2_u4_u4_n143 ) , .A( u2_u4_u4_n174 ) , .B1( u2_u4_u4_n184 ) );
  AOI21_X1 u2_u4_u4_U15 (.B2( u2_u4_u4_n158 ) , .B1( u2_u4_u4_n159 ) , .ZN( u2_u4_u4_n163 ) , .A( u2_u4_u4_n174 ) );
  AOI21_X1 u2_u4_u4_U16 (.A( u2_u4_u4_n153 ) , .B2( u2_u4_u4_n154 ) , .B1( u2_u4_u4_n155 ) , .ZN( u2_u4_u4_n165 ) );
  AOI21_X1 u2_u4_u4_U17 (.A( u2_u4_u4_n156 ) , .B2( u2_u4_u4_n157 ) , .ZN( u2_u4_u4_n164 ) , .B1( u2_u4_u4_n184 ) );
  INV_X1 u2_u4_u4_U18 (.A( u2_u4_u4_n138 ) , .ZN( u2_u4_u4_n170 ) );
  AND2_X1 u2_u4_u4_U19 (.A2( u2_u4_u4_n120 ) , .ZN( u2_u4_u4_n155 ) , .A1( u2_u4_u4_n160 ) );
  INV_X1 u2_u4_u4_U20 (.A( u2_u4_u4_n156 ) , .ZN( u2_u4_u4_n175 ) );
  NAND2_X1 u2_u4_u4_U21 (.A2( u2_u4_u4_n118 ) , .ZN( u2_u4_u4_n131 ) , .A1( u2_u4_u4_n147 ) );
  NAND2_X1 u2_u4_u4_U22 (.A1( u2_u4_u4_n119 ) , .A2( u2_u4_u4_n120 ) , .ZN( u2_u4_u4_n130 ) );
  NAND2_X1 u2_u4_u4_U23 (.ZN( u2_u4_u4_n117 ) , .A2( u2_u4_u4_n118 ) , .A1( u2_u4_u4_n148 ) );
  NAND2_X1 u2_u4_u4_U24 (.ZN( u2_u4_u4_n129 ) , .A1( u2_u4_u4_n134 ) , .A2( u2_u4_u4_n148 ) );
  AND3_X1 u2_u4_u4_U25 (.A1( u2_u4_u4_n119 ) , .A2( u2_u4_u4_n143 ) , .A3( u2_u4_u4_n154 ) , .ZN( u2_u4_u4_n161 ) );
  AND2_X1 u2_u4_u4_U26 (.A1( u2_u4_u4_n145 ) , .A2( u2_u4_u4_n147 ) , .ZN( u2_u4_u4_n159 ) );
  OR3_X1 u2_u4_u4_U27 (.A3( u2_u4_u4_n114 ) , .A2( u2_u4_u4_n115 ) , .A1( u2_u4_u4_n116 ) , .ZN( u2_u4_u4_n136 ) );
  AOI21_X1 u2_u4_u4_U28 (.A( u2_u4_u4_n113 ) , .ZN( u2_u4_u4_n116 ) , .B2( u2_u4_u4_n173 ) , .B1( u2_u4_u4_n174 ) );
  AOI21_X1 u2_u4_u4_U29 (.ZN( u2_u4_u4_n115 ) , .B2( u2_u4_u4_n145 ) , .B1( u2_u4_u4_n146 ) , .A( u2_u4_u4_n156 ) );
  NOR2_X1 u2_u4_u4_U3 (.ZN( u2_u4_u4_n121 ) , .A1( u2_u4_u4_n181 ) , .A2( u2_u4_u4_n182 ) );
  OAI22_X1 u2_u4_u4_U30 (.ZN( u2_u4_u4_n114 ) , .A2( u2_u4_u4_n121 ) , .B1( u2_u4_u4_n160 ) , .B2( u2_u4_u4_n170 ) , .A1( u2_u4_u4_n171 ) );
  INV_X1 u2_u4_u4_U31 (.A( u2_u4_u4_n158 ) , .ZN( u2_u4_u4_n182 ) );
  INV_X1 u2_u4_u4_U32 (.ZN( u2_u4_u4_n181 ) , .A( u2_u4_u4_n96 ) );
  INV_X1 u2_u4_u4_U33 (.A( u2_u4_u4_n144 ) , .ZN( u2_u4_u4_n179 ) );
  INV_X1 u2_u4_u4_U34 (.A( u2_u4_u4_n157 ) , .ZN( u2_u4_u4_n178 ) );
  NAND2_X1 u2_u4_u4_U35 (.A2( u2_u4_u4_n154 ) , .A1( u2_u4_u4_n96 ) , .ZN( u2_u4_u4_n97 ) );
  INV_X1 u2_u4_u4_U36 (.ZN( u2_u4_u4_n186 ) , .A( u2_u4_u4_n95 ) );
  OAI221_X1 u2_u4_u4_U37 (.C1( u2_u4_u4_n134 ) , .B1( u2_u4_u4_n158 ) , .B2( u2_u4_u4_n171 ) , .C2( u2_u4_u4_n173 ) , .A( u2_u4_u4_n94 ) , .ZN( u2_u4_u4_n95 ) );
  AOI222_X1 u2_u4_u4_U38 (.B2( u2_u4_u4_n132 ) , .A1( u2_u4_u4_n138 ) , .C2( u2_u4_u4_n175 ) , .A2( u2_u4_u4_n179 ) , .C1( u2_u4_u4_n181 ) , .B1( u2_u4_u4_n185 ) , .ZN( u2_u4_u4_n94 ) );
  INV_X1 u2_u4_u4_U39 (.A( u2_u4_u4_n113 ) , .ZN( u2_u4_u4_n185 ) );
  INV_X1 u2_u4_u4_U4 (.A( u2_u4_u4_n117 ) , .ZN( u2_u4_u4_n184 ) );
  INV_X1 u2_u4_u4_U40 (.A( u2_u4_u4_n143 ) , .ZN( u2_u4_u4_n183 ) );
  NOR2_X1 u2_u4_u4_U41 (.ZN( u2_u4_u4_n138 ) , .A1( u2_u4_u4_n168 ) , .A2( u2_u4_u4_n169 ) );
  NOR2_X1 u2_u4_u4_U42 (.A1( u2_u4_u4_n150 ) , .A2( u2_u4_u4_n152 ) , .ZN( u2_u4_u4_n153 ) );
  NOR2_X1 u2_u4_u4_U43 (.A2( u2_u4_u4_n128 ) , .A1( u2_u4_u4_n138 ) , .ZN( u2_u4_u4_n156 ) );
  AOI22_X1 u2_u4_u4_U44 (.B2( u2_u4_u4_n122 ) , .A1( u2_u4_u4_n123 ) , .ZN( u2_u4_u4_n124 ) , .B1( u2_u4_u4_n128 ) , .A2( u2_u4_u4_n172 ) );
  INV_X1 u2_u4_u4_U45 (.A( u2_u4_u4_n153 ) , .ZN( u2_u4_u4_n172 ) );
  NAND2_X1 u2_u4_u4_U46 (.A2( u2_u4_u4_n120 ) , .ZN( u2_u4_u4_n123 ) , .A1( u2_u4_u4_n161 ) );
  AOI22_X1 u2_u4_u4_U47 (.B2( u2_u4_u4_n132 ) , .A2( u2_u4_u4_n133 ) , .ZN( u2_u4_u4_n140 ) , .A1( u2_u4_u4_n150 ) , .B1( u2_u4_u4_n179 ) );
  NAND2_X1 u2_u4_u4_U48 (.ZN( u2_u4_u4_n133 ) , .A2( u2_u4_u4_n146 ) , .A1( u2_u4_u4_n154 ) );
  NAND2_X1 u2_u4_u4_U49 (.A1( u2_u4_u4_n103 ) , .ZN( u2_u4_u4_n154 ) , .A2( u2_u4_u4_n98 ) );
  NOR4_X1 u2_u4_u4_U5 (.A4( u2_u4_u4_n106 ) , .A3( u2_u4_u4_n107 ) , .A2( u2_u4_u4_n108 ) , .A1( u2_u4_u4_n109 ) , .ZN( u2_u4_u4_n110 ) );
  NAND2_X1 u2_u4_u4_U50 (.A1( u2_u4_u4_n101 ) , .ZN( u2_u4_u4_n158 ) , .A2( u2_u4_u4_n99 ) );
  AOI21_X1 u2_u4_u4_U51 (.ZN( u2_u4_u4_n127 ) , .A( u2_u4_u4_n136 ) , .B2( u2_u4_u4_n150 ) , .B1( u2_u4_u4_n180 ) );
  INV_X1 u2_u4_u4_U52 (.A( u2_u4_u4_n160 ) , .ZN( u2_u4_u4_n180 ) );
  NAND2_X1 u2_u4_u4_U53 (.A2( u2_u4_u4_n104 ) , .A1( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n146 ) );
  NAND2_X1 u2_u4_u4_U54 (.A2( u2_u4_u4_n101 ) , .A1( u2_u4_u4_n102 ) , .ZN( u2_u4_u4_n160 ) );
  NAND2_X1 u2_u4_u4_U55 (.ZN( u2_u4_u4_n134 ) , .A1( u2_u4_u4_n98 ) , .A2( u2_u4_u4_n99 ) );
  NAND2_X1 u2_u4_u4_U56 (.A1( u2_u4_u4_n103 ) , .A2( u2_u4_u4_n104 ) , .ZN( u2_u4_u4_n143 ) );
  NAND2_X1 u2_u4_u4_U57 (.A2( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n145 ) , .A1( u2_u4_u4_n98 ) );
  NAND2_X1 u2_u4_u4_U58 (.A1( u2_u4_u4_n100 ) , .A2( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n120 ) );
  NAND2_X1 u2_u4_u4_U59 (.A1( u2_u4_u4_n102 ) , .A2( u2_u4_u4_n104 ) , .ZN( u2_u4_u4_n148 ) );
  AOI21_X1 u2_u4_u4_U6 (.ZN( u2_u4_u4_n106 ) , .B2( u2_u4_u4_n146 ) , .B1( u2_u4_u4_n158 ) , .A( u2_u4_u4_n170 ) );
  NAND2_X1 u2_u4_u4_U60 (.A2( u2_u4_u4_n100 ) , .A1( u2_u4_u4_n103 ) , .ZN( u2_u4_u4_n157 ) );
  INV_X1 u2_u4_u4_U61 (.A( u2_u4_u4_n150 ) , .ZN( u2_u4_u4_n173 ) );
  INV_X1 u2_u4_u4_U62 (.A( u2_u4_u4_n152 ) , .ZN( u2_u4_u4_n171 ) );
  NAND2_X1 u2_u4_u4_U63 (.A1( u2_u4_u4_n100 ) , .ZN( u2_u4_u4_n118 ) , .A2( u2_u4_u4_n99 ) );
  NAND2_X1 u2_u4_u4_U64 (.A2( u2_u4_u4_n100 ) , .A1( u2_u4_u4_n102 ) , .ZN( u2_u4_u4_n144 ) );
  NAND2_X1 u2_u4_u4_U65 (.A2( u2_u4_u4_n101 ) , .A1( u2_u4_u4_n105 ) , .ZN( u2_u4_u4_n96 ) );
  INV_X1 u2_u4_u4_U66 (.A( u2_u4_u4_n128 ) , .ZN( u2_u4_u4_n174 ) );
  NAND2_X1 u2_u4_u4_U67 (.A2( u2_u4_u4_n102 ) , .ZN( u2_u4_u4_n119 ) , .A1( u2_u4_u4_n98 ) );
  NAND2_X1 u2_u4_u4_U68 (.A2( u2_u4_u4_n101 ) , .A1( u2_u4_u4_n103 ) , .ZN( u2_u4_u4_n147 ) );
  NAND2_X1 u2_u4_u4_U69 (.A2( u2_u4_u4_n104 ) , .ZN( u2_u4_u4_n113 ) , .A1( u2_u4_u4_n99 ) );
  AOI21_X1 u2_u4_u4_U7 (.ZN( u2_u4_u4_n108 ) , .B2( u2_u4_u4_n134 ) , .B1( u2_u4_u4_n155 ) , .A( u2_u4_u4_n156 ) );
  NOR2_X1 u2_u4_u4_U70 (.A2( u2_u4_X_28 ) , .ZN( u2_u4_u4_n150 ) , .A1( u2_u4_u4_n168 ) );
  NOR2_X1 u2_u4_u4_U71 (.A2( u2_u4_X_29 ) , .ZN( u2_u4_u4_n152 ) , .A1( u2_u4_u4_n169 ) );
  NOR2_X1 u2_u4_u4_U72 (.A2( u2_u4_X_30 ) , .ZN( u2_u4_u4_n105 ) , .A1( u2_u4_u4_n176 ) );
  NOR2_X1 u2_u4_u4_U73 (.A2( u2_u4_X_26 ) , .ZN( u2_u4_u4_n100 ) , .A1( u2_u4_u4_n177 ) );
  NOR2_X1 u2_u4_u4_U74 (.A2( u2_u4_X_28 ) , .A1( u2_u4_X_29 ) , .ZN( u2_u4_u4_n128 ) );
  NOR2_X1 u2_u4_u4_U75 (.A2( u2_u4_X_27 ) , .A1( u2_u4_X_30 ) , .ZN( u2_u4_u4_n102 ) );
  NOR2_X1 u2_u4_u4_U76 (.A2( u2_u4_X_25 ) , .A1( u2_u4_X_26 ) , .ZN( u2_u4_u4_n98 ) );
  AND2_X1 u2_u4_u4_U77 (.A2( u2_u4_X_25 ) , .A1( u2_u4_X_26 ) , .ZN( u2_u4_u4_n104 ) );
  AND2_X1 u2_u4_u4_U78 (.A1( u2_u4_X_30 ) , .A2( u2_u4_u4_n176 ) , .ZN( u2_u4_u4_n99 ) );
  AND2_X1 u2_u4_u4_U79 (.A1( u2_u4_X_26 ) , .ZN( u2_u4_u4_n101 ) , .A2( u2_u4_u4_n177 ) );
  AOI21_X1 u2_u4_u4_U8 (.ZN( u2_u4_u4_n109 ) , .A( u2_u4_u4_n153 ) , .B1( u2_u4_u4_n159 ) , .B2( u2_u4_u4_n184 ) );
  AND2_X1 u2_u4_u4_U80 (.A1( u2_u4_X_27 ) , .A2( u2_u4_X_30 ) , .ZN( u2_u4_u4_n103 ) );
  INV_X1 u2_u4_u4_U81 (.A( u2_u4_X_28 ) , .ZN( u2_u4_u4_n169 ) );
  INV_X1 u2_u4_u4_U82 (.A( u2_u4_X_29 ) , .ZN( u2_u4_u4_n168 ) );
  INV_X1 u2_u4_u4_U83 (.A( u2_u4_X_25 ) , .ZN( u2_u4_u4_n177 ) );
  INV_X1 u2_u4_u4_U84 (.A( u2_u4_X_27 ) , .ZN( u2_u4_u4_n176 ) );
  NAND4_X1 u2_u4_u4_U85 (.ZN( u2_out4_25 ) , .A4( u2_u4_u4_n139 ) , .A3( u2_u4_u4_n140 ) , .A2( u2_u4_u4_n141 ) , .A1( u2_u4_u4_n142 ) );
  OAI21_X1 u2_u4_u4_U86 (.B2( u2_u4_u4_n131 ) , .ZN( u2_u4_u4_n141 ) , .A( u2_u4_u4_n175 ) , .B1( u2_u4_u4_n183 ) );
  OAI21_X1 u2_u4_u4_U87 (.A( u2_u4_u4_n128 ) , .B2( u2_u4_u4_n129 ) , .B1( u2_u4_u4_n130 ) , .ZN( u2_u4_u4_n142 ) );
  NAND4_X1 u2_u4_u4_U88 (.ZN( u2_out4_14 ) , .A4( u2_u4_u4_n124 ) , .A3( u2_u4_u4_n125 ) , .A2( u2_u4_u4_n126 ) , .A1( u2_u4_u4_n127 ) );
  AOI22_X1 u2_u4_u4_U89 (.B2( u2_u4_u4_n117 ) , .ZN( u2_u4_u4_n126 ) , .A1( u2_u4_u4_n129 ) , .B1( u2_u4_u4_n152 ) , .A2( u2_u4_u4_n175 ) );
  AOI211_X1 u2_u4_u4_U9 (.B( u2_u4_u4_n136 ) , .A( u2_u4_u4_n137 ) , .C2( u2_u4_u4_n138 ) , .ZN( u2_u4_u4_n139 ) , .C1( u2_u4_u4_n182 ) );
  AOI22_X1 u2_u4_u4_U90 (.ZN( u2_u4_u4_n125 ) , .B2( u2_u4_u4_n131 ) , .A2( u2_u4_u4_n132 ) , .B1( u2_u4_u4_n138 ) , .A1( u2_u4_u4_n178 ) );
  NAND4_X1 u2_u4_u4_U91 (.ZN( u2_out4_8 ) , .A4( u2_u4_u4_n110 ) , .A3( u2_u4_u4_n111 ) , .A2( u2_u4_u4_n112 ) , .A1( u2_u4_u4_n186 ) );
  NAND2_X1 u2_u4_u4_U92 (.ZN( u2_u4_u4_n112 ) , .A2( u2_u4_u4_n130 ) , .A1( u2_u4_u4_n150 ) );
  AOI22_X1 u2_u4_u4_U93 (.ZN( u2_u4_u4_n111 ) , .B2( u2_u4_u4_n132 ) , .A1( u2_u4_u4_n152 ) , .B1( u2_u4_u4_n178 ) , .A2( u2_u4_u4_n97 ) );
  AOI22_X1 u2_u4_u4_U94 (.B2( u2_u4_u4_n149 ) , .B1( u2_u4_u4_n150 ) , .A2( u2_u4_u4_n151 ) , .A1( u2_u4_u4_n152 ) , .ZN( u2_u4_u4_n167 ) );
  NOR4_X1 u2_u4_u4_U95 (.A4( u2_u4_u4_n162 ) , .A3( u2_u4_u4_n163 ) , .A2( u2_u4_u4_n164 ) , .A1( u2_u4_u4_n165 ) , .ZN( u2_u4_u4_n166 ) );
  NAND3_X1 u2_u4_u4_U96 (.ZN( u2_out4_3 ) , .A3( u2_u4_u4_n166 ) , .A1( u2_u4_u4_n167 ) , .A2( u2_u4_u4_n186 ) );
  NAND3_X1 u2_u4_u4_U97 (.A3( u2_u4_u4_n146 ) , .A2( u2_u4_u4_n147 ) , .A1( u2_u4_u4_n148 ) , .ZN( u2_u4_u4_n149 ) );
  NAND3_X1 u2_u4_u4_U98 (.A3( u2_u4_u4_n143 ) , .A2( u2_u4_u4_n144 ) , .A1( u2_u4_u4_n145 ) , .ZN( u2_u4_u4_n151 ) );
  NAND3_X1 u2_u4_u4_U99 (.A3( u2_u4_u4_n121 ) , .ZN( u2_u4_u4_n122 ) , .A2( u2_u4_u4_n144 ) , .A1( u2_u4_u4_n154 ) );
  XOR2_X1 u2_u7_U16 (.B( u2_K8_3 ) , .A( u2_R6_2 ) , .Z( u2_u7_X_3 ) );
  XOR2_X1 u2_u7_U27 (.B( u2_K8_2 ) , .A( u2_R6_1 ) , .Z( u2_u7_X_2 ) );
  XOR2_X1 u2_u7_U38 (.B( u2_K8_1 ) , .A( u2_R6_32 ) , .Z( u2_u7_X_1 ) );
  XOR2_X1 u2_u7_U4 (.B( u2_K8_6 ) , .A( u2_R6_5 ) , .Z( u2_u7_X_6 ) );
  XOR2_X1 u2_u7_U40 (.B( u2_K8_18 ) , .A( u2_R6_13 ) , .Z( u2_u7_X_18 ) );
  XOR2_X1 u2_u7_U41 (.B( u2_K8_17 ) , .A( u2_R6_12 ) , .Z( u2_u7_X_17 ) );
  XOR2_X1 u2_u7_U42 (.B( u2_K8_16 ) , .A( u2_R6_11 ) , .Z( u2_u7_X_16 ) );
  XOR2_X1 u2_u7_U43 (.B( u2_K8_15 ) , .A( u2_R6_10 ) , .Z( u2_u7_X_15 ) );
  XOR2_X1 u2_u7_U44 (.B( u2_K8_14 ) , .A( u2_R6_9 ) , .Z( u2_u7_X_14 ) );
  XOR2_X1 u2_u7_U45 (.B( u2_K8_13 ) , .A( u2_R6_8 ) , .Z( u2_u7_X_13 ) );
  XOR2_X1 u2_u7_U5 (.B( u2_K8_5 ) , .A( u2_R6_4 ) , .Z( u2_u7_X_5 ) );
  XOR2_X1 u2_u7_U6 (.B( u2_K8_4 ) , .A( u2_R6_3 ) , .Z( u2_u7_X_4 ) );
  AND3_X1 u2_u7_u0_U10 (.A2( u2_u7_u0_n112 ) , .ZN( u2_u7_u0_n127 ) , .A3( u2_u7_u0_n130 ) , .A1( u2_u7_u0_n148 ) );
  NAND2_X1 u2_u7_u0_U11 (.ZN( u2_u7_u0_n113 ) , .A1( u2_u7_u0_n139 ) , .A2( u2_u7_u0_n149 ) );
  AND2_X1 u2_u7_u0_U12 (.ZN( u2_u7_u0_n107 ) , .A1( u2_u7_u0_n130 ) , .A2( u2_u7_u0_n140 ) );
  AND2_X1 u2_u7_u0_U13 (.A2( u2_u7_u0_n129 ) , .A1( u2_u7_u0_n130 ) , .ZN( u2_u7_u0_n151 ) );
  AND2_X1 u2_u7_u0_U14 (.A1( u2_u7_u0_n108 ) , .A2( u2_u7_u0_n125 ) , .ZN( u2_u7_u0_n145 ) );
  INV_X1 u2_u7_u0_U15 (.A( u2_u7_u0_n143 ) , .ZN( u2_u7_u0_n173 ) );
  NOR2_X1 u2_u7_u0_U16 (.A2( u2_u7_u0_n136 ) , .ZN( u2_u7_u0_n147 ) , .A1( u2_u7_u0_n160 ) );
  INV_X1 u2_u7_u0_U17 (.ZN( u2_u7_u0_n172 ) , .A( u2_u7_u0_n88 ) );
  OAI222_X1 u2_u7_u0_U18 (.C1( u2_u7_u0_n108 ) , .A1( u2_u7_u0_n125 ) , .B2( u2_u7_u0_n128 ) , .B1( u2_u7_u0_n144 ) , .A2( u2_u7_u0_n158 ) , .C2( u2_u7_u0_n161 ) , .ZN( u2_u7_u0_n88 ) );
  NOR2_X1 u2_u7_u0_U19 (.A1( u2_u7_u0_n163 ) , .A2( u2_u7_u0_n164 ) , .ZN( u2_u7_u0_n95 ) );
  OAI22_X1 u2_u7_u0_U20 (.B1( u2_u7_u0_n125 ) , .ZN( u2_u7_u0_n126 ) , .A1( u2_u7_u0_n138 ) , .A2( u2_u7_u0_n146 ) , .B2( u2_u7_u0_n147 ) );
  OAI22_X1 u2_u7_u0_U21 (.B1( u2_u7_u0_n131 ) , .A1( u2_u7_u0_n144 ) , .B2( u2_u7_u0_n147 ) , .A2( u2_u7_u0_n90 ) , .ZN( u2_u7_u0_n91 ) );
  AND3_X1 u2_u7_u0_U22 (.A3( u2_u7_u0_n121 ) , .A2( u2_u7_u0_n125 ) , .A1( u2_u7_u0_n148 ) , .ZN( u2_u7_u0_n90 ) );
  INV_X1 u2_u7_u0_U23 (.A( u2_u7_u0_n136 ) , .ZN( u2_u7_u0_n161 ) );
  AOI22_X1 u2_u7_u0_U24 (.B2( u2_u7_u0_n109 ) , .A2( u2_u7_u0_n110 ) , .ZN( u2_u7_u0_n111 ) , .B1( u2_u7_u0_n118 ) , .A1( u2_u7_u0_n160 ) );
  INV_X1 u2_u7_u0_U25 (.A( u2_u7_u0_n118 ) , .ZN( u2_u7_u0_n158 ) );
  AOI21_X1 u2_u7_u0_U26 (.ZN( u2_u7_u0_n104 ) , .B1( u2_u7_u0_n107 ) , .B2( u2_u7_u0_n141 ) , .A( u2_u7_u0_n144 ) );
  AOI21_X1 u2_u7_u0_U27 (.B1( u2_u7_u0_n127 ) , .B2( u2_u7_u0_n129 ) , .A( u2_u7_u0_n138 ) , .ZN( u2_u7_u0_n96 ) );
  AOI21_X1 u2_u7_u0_U28 (.ZN( u2_u7_u0_n116 ) , .B2( u2_u7_u0_n142 ) , .A( u2_u7_u0_n144 ) , .B1( u2_u7_u0_n166 ) );
  INV_X1 u2_u7_u0_U29 (.ZN( u2_u7_u0_n171 ) , .A( u2_u7_u0_n99 ) );
  INV_X1 u2_u7_u0_U3 (.A( u2_u7_u0_n113 ) , .ZN( u2_u7_u0_n166 ) );
  OAI211_X1 u2_u7_u0_U30 (.C2( u2_u7_u0_n140 ) , .C1( u2_u7_u0_n161 ) , .A( u2_u7_u0_n169 ) , .B( u2_u7_u0_n98 ) , .ZN( u2_u7_u0_n99 ) );
  INV_X1 u2_u7_u0_U31 (.ZN( u2_u7_u0_n169 ) , .A( u2_u7_u0_n91 ) );
  AOI211_X1 u2_u7_u0_U32 (.C1( u2_u7_u0_n118 ) , .A( u2_u7_u0_n123 ) , .B( u2_u7_u0_n96 ) , .C2( u2_u7_u0_n97 ) , .ZN( u2_u7_u0_n98 ) );
  NOR2_X1 u2_u7_u0_U33 (.A1( u2_u7_u0_n120 ) , .ZN( u2_u7_u0_n143 ) , .A2( u2_u7_u0_n167 ) );
  OAI221_X1 u2_u7_u0_U34 (.C1( u2_u7_u0_n112 ) , .ZN( u2_u7_u0_n120 ) , .B1( u2_u7_u0_n138 ) , .B2( u2_u7_u0_n141 ) , .C2( u2_u7_u0_n147 ) , .A( u2_u7_u0_n172 ) );
  AOI211_X1 u2_u7_u0_U35 (.B( u2_u7_u0_n115 ) , .A( u2_u7_u0_n116 ) , .C2( u2_u7_u0_n117 ) , .C1( u2_u7_u0_n118 ) , .ZN( u2_u7_u0_n119 ) );
  NAND2_X1 u2_u7_u0_U36 (.A1( u2_u7_u0_n101 ) , .A2( u2_u7_u0_n102 ) , .ZN( u2_u7_u0_n150 ) );
  INV_X1 u2_u7_u0_U37 (.A( u2_u7_u0_n138 ) , .ZN( u2_u7_u0_n160 ) );
  NAND2_X1 u2_u7_u0_U38 (.A1( u2_u7_u0_n102 ) , .ZN( u2_u7_u0_n128 ) , .A2( u2_u7_u0_n95 ) );
  NAND2_X1 u2_u7_u0_U39 (.ZN( u2_u7_u0_n148 ) , .A1( u2_u7_u0_n93 ) , .A2( u2_u7_u0_n95 ) );
  AOI21_X1 u2_u7_u0_U4 (.B1( u2_u7_u0_n114 ) , .ZN( u2_u7_u0_n115 ) , .B2( u2_u7_u0_n129 ) , .A( u2_u7_u0_n161 ) );
  NAND2_X1 u2_u7_u0_U40 (.A2( u2_u7_u0_n102 ) , .A1( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n149 ) );
  NAND2_X1 u2_u7_u0_U41 (.A2( u2_u7_u0_n102 ) , .ZN( u2_u7_u0_n114 ) , .A1( u2_u7_u0_n92 ) );
  NAND2_X1 u2_u7_u0_U42 (.A2( u2_u7_u0_n101 ) , .ZN( u2_u7_u0_n121 ) , .A1( u2_u7_u0_n93 ) );
  NAND2_X1 u2_u7_u0_U43 (.ZN( u2_u7_u0_n112 ) , .A2( u2_u7_u0_n92 ) , .A1( u2_u7_u0_n93 ) );
  AOI21_X1 u2_u7_u0_U44 (.B1( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n132 ) , .A( u2_u7_u0_n165 ) , .B2( u2_u7_u0_n93 ) );
  INV_X1 u2_u7_u0_U45 (.A( u2_u7_u0_n142 ) , .ZN( u2_u7_u0_n165 ) );
  OR3_X1 u2_u7_u0_U46 (.A3( u2_u7_u0_n152 ) , .A2( u2_u7_u0_n153 ) , .A1( u2_u7_u0_n154 ) , .ZN( u2_u7_u0_n155 ) );
  AOI21_X1 u2_u7_u0_U47 (.A( u2_u7_u0_n144 ) , .B2( u2_u7_u0_n145 ) , .B1( u2_u7_u0_n146 ) , .ZN( u2_u7_u0_n154 ) );
  AOI21_X1 u2_u7_u0_U48 (.B2( u2_u7_u0_n150 ) , .B1( u2_u7_u0_n151 ) , .ZN( u2_u7_u0_n152 ) , .A( u2_u7_u0_n158 ) );
  AOI21_X1 u2_u7_u0_U49 (.A( u2_u7_u0_n147 ) , .B2( u2_u7_u0_n148 ) , .B1( u2_u7_u0_n149 ) , .ZN( u2_u7_u0_n153 ) );
  AOI21_X1 u2_u7_u0_U5 (.B2( u2_u7_u0_n131 ) , .ZN( u2_u7_u0_n134 ) , .B1( u2_u7_u0_n151 ) , .A( u2_u7_u0_n158 ) );
  NOR2_X1 u2_u7_u0_U50 (.A2( u2_u7_X_4 ) , .A1( u2_u7_X_5 ) , .ZN( u2_u7_u0_n118 ) );
  NAND2_X1 u2_u7_u0_U51 (.A2( u2_u7_X_4 ) , .A1( u2_u7_X_5 ) , .ZN( u2_u7_u0_n144 ) );
  NOR2_X1 u2_u7_u0_U52 (.A2( u2_u7_X_1 ) , .A1( u2_u7_X_2 ) , .ZN( u2_u7_u0_n92 ) );
  NOR2_X1 u2_u7_u0_U53 (.A2( u2_u7_X_1 ) , .ZN( u2_u7_u0_n101 ) , .A1( u2_u7_u0_n163 ) );
  NOR2_X1 u2_u7_u0_U54 (.A2( u2_u7_X_2 ) , .ZN( u2_u7_u0_n103 ) , .A1( u2_u7_u0_n164 ) );
  NOR2_X1 u2_u7_u0_U55 (.A2( u2_u7_X_5 ) , .ZN( u2_u7_u0_n136 ) , .A1( u2_u7_u0_n159 ) );
  NAND2_X1 u2_u7_u0_U56 (.A1( u2_u7_X_5 ) , .ZN( u2_u7_u0_n138 ) , .A2( u2_u7_u0_n159 ) );
  AND2_X1 u2_u7_u0_U57 (.A2( u2_u7_X_3 ) , .A1( u2_u7_X_6 ) , .ZN( u2_u7_u0_n102 ) );
  AND2_X1 u2_u7_u0_U58 (.A1( u2_u7_X_6 ) , .A2( u2_u7_u0_n162 ) , .ZN( u2_u7_u0_n93 ) );
  INV_X1 u2_u7_u0_U59 (.A( u2_u7_X_4 ) , .ZN( u2_u7_u0_n159 ) );
  NOR2_X1 u2_u7_u0_U6 (.A1( u2_u7_u0_n108 ) , .ZN( u2_u7_u0_n123 ) , .A2( u2_u7_u0_n158 ) );
  INV_X1 u2_u7_u0_U60 (.A( u2_u7_X_1 ) , .ZN( u2_u7_u0_n164 ) );
  INV_X1 u2_u7_u0_U61 (.A( u2_u7_X_2 ) , .ZN( u2_u7_u0_n163 ) );
  INV_X1 u2_u7_u0_U62 (.A( u2_u7_u0_n126 ) , .ZN( u2_u7_u0_n168 ) );
  AOI211_X1 u2_u7_u0_U63 (.B( u2_u7_u0_n133 ) , .A( u2_u7_u0_n134 ) , .C2( u2_u7_u0_n135 ) , .C1( u2_u7_u0_n136 ) , .ZN( u2_u7_u0_n137 ) );
  OR4_X1 u2_u7_u0_U64 (.ZN( u2_out7_17 ) , .A4( u2_u7_u0_n122 ) , .A2( u2_u7_u0_n123 ) , .A1( u2_u7_u0_n124 ) , .A3( u2_u7_u0_n170 ) );
  AOI21_X1 u2_u7_u0_U65 (.B2( u2_u7_u0_n107 ) , .ZN( u2_u7_u0_n124 ) , .B1( u2_u7_u0_n128 ) , .A( u2_u7_u0_n161 ) );
  INV_X1 u2_u7_u0_U66 (.A( u2_u7_u0_n111 ) , .ZN( u2_u7_u0_n170 ) );
  OR4_X1 u2_u7_u0_U67 (.ZN( u2_out7_31 ) , .A4( u2_u7_u0_n155 ) , .A2( u2_u7_u0_n156 ) , .A1( u2_u7_u0_n157 ) , .A3( u2_u7_u0_n173 ) );
  AOI21_X1 u2_u7_u0_U68 (.A( u2_u7_u0_n138 ) , .B2( u2_u7_u0_n139 ) , .B1( u2_u7_u0_n140 ) , .ZN( u2_u7_u0_n157 ) );
  AOI21_X1 u2_u7_u0_U69 (.B2( u2_u7_u0_n141 ) , .B1( u2_u7_u0_n142 ) , .ZN( u2_u7_u0_n156 ) , .A( u2_u7_u0_n161 ) );
  OAI21_X1 u2_u7_u0_U7 (.B1( u2_u7_u0_n150 ) , .B2( u2_u7_u0_n158 ) , .A( u2_u7_u0_n172 ) , .ZN( u2_u7_u0_n89 ) );
  INV_X1 u2_u7_u0_U70 (.ZN( u2_u7_u0_n174 ) , .A( u2_u7_u0_n89 ) );
  AOI211_X1 u2_u7_u0_U71 (.B( u2_u7_u0_n104 ) , .A( u2_u7_u0_n105 ) , .ZN( u2_u7_u0_n106 ) , .C2( u2_u7_u0_n113 ) , .C1( u2_u7_u0_n160 ) );
  NAND2_X1 u2_u7_u0_U72 (.A2( u2_u7_u0_n100 ) , .A1( u2_u7_u0_n101 ) , .ZN( u2_u7_u0_n139 ) );
  NAND2_X1 u2_u7_u0_U73 (.A1( u2_u7_u0_n100 ) , .A2( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n125 ) );
  NAND2_X1 u2_u7_u0_U74 (.A1( u2_u7_u0_n100 ) , .ZN( u2_u7_u0_n129 ) , .A2( u2_u7_u0_n95 ) );
  NAND2_X1 u2_u7_u0_U75 (.A2( u2_u7_u0_n100 ) , .ZN( u2_u7_u0_n131 ) , .A1( u2_u7_u0_n92 ) );
  OAI221_X1 u2_u7_u0_U76 (.C1( u2_u7_u0_n121 ) , .ZN( u2_u7_u0_n122 ) , .B2( u2_u7_u0_n127 ) , .A( u2_u7_u0_n143 ) , .B1( u2_u7_u0_n144 ) , .C2( u2_u7_u0_n147 ) );
  NOR2_X1 u2_u7_u0_U77 (.A2( u2_u7_X_6 ) , .ZN( u2_u7_u0_n100 ) , .A1( u2_u7_u0_n162 ) );
  AOI21_X1 u2_u7_u0_U78 (.B1( u2_u7_u0_n132 ) , .ZN( u2_u7_u0_n133 ) , .A( u2_u7_u0_n144 ) , .B2( u2_u7_u0_n166 ) );
  OAI22_X1 u2_u7_u0_U79 (.ZN( u2_u7_u0_n105 ) , .A2( u2_u7_u0_n132 ) , .B1( u2_u7_u0_n146 ) , .A1( u2_u7_u0_n147 ) , .B2( u2_u7_u0_n161 ) );
  AND2_X1 u2_u7_u0_U8 (.A1( u2_u7_u0_n114 ) , .A2( u2_u7_u0_n121 ) , .ZN( u2_u7_u0_n146 ) );
  NAND2_X1 u2_u7_u0_U80 (.ZN( u2_u7_u0_n110 ) , .A2( u2_u7_u0_n132 ) , .A1( u2_u7_u0_n145 ) );
  INV_X1 u2_u7_u0_U81 (.A( u2_u7_u0_n119 ) , .ZN( u2_u7_u0_n167 ) );
  NAND2_X1 u2_u7_u0_U82 (.A2( u2_u7_u0_n103 ) , .ZN( u2_u7_u0_n140 ) , .A1( u2_u7_u0_n94 ) );
  NAND2_X1 u2_u7_u0_U83 (.A1( u2_u7_u0_n101 ) , .ZN( u2_u7_u0_n130 ) , .A2( u2_u7_u0_n94 ) );
  NAND2_X1 u2_u7_u0_U84 (.ZN( u2_u7_u0_n108 ) , .A1( u2_u7_u0_n92 ) , .A2( u2_u7_u0_n94 ) );
  NAND2_X1 u2_u7_u0_U85 (.ZN( u2_u7_u0_n142 ) , .A1( u2_u7_u0_n94 ) , .A2( u2_u7_u0_n95 ) );
  INV_X1 u2_u7_u0_U86 (.A( u2_u7_X_3 ) , .ZN( u2_u7_u0_n162 ) );
  NOR2_X1 u2_u7_u0_U87 (.A2( u2_u7_X_3 ) , .A1( u2_u7_X_6 ) , .ZN( u2_u7_u0_n94 ) );
  NAND3_X1 u2_u7_u0_U88 (.ZN( u2_out7_23 ) , .A3( u2_u7_u0_n137 ) , .A1( u2_u7_u0_n168 ) , .A2( u2_u7_u0_n171 ) );
  NAND3_X1 u2_u7_u0_U89 (.A3( u2_u7_u0_n127 ) , .A2( u2_u7_u0_n128 ) , .ZN( u2_u7_u0_n135 ) , .A1( u2_u7_u0_n150 ) );
  AND2_X1 u2_u7_u0_U9 (.A1( u2_u7_u0_n131 ) , .ZN( u2_u7_u0_n141 ) , .A2( u2_u7_u0_n150 ) );
  NAND3_X1 u2_u7_u0_U90 (.ZN( u2_u7_u0_n117 ) , .A3( u2_u7_u0_n132 ) , .A2( u2_u7_u0_n139 ) , .A1( u2_u7_u0_n148 ) );
  NAND3_X1 u2_u7_u0_U91 (.ZN( u2_u7_u0_n109 ) , .A2( u2_u7_u0_n114 ) , .A3( u2_u7_u0_n140 ) , .A1( u2_u7_u0_n149 ) );
  NAND3_X1 u2_u7_u0_U92 (.ZN( u2_out7_9 ) , .A3( u2_u7_u0_n106 ) , .A2( u2_u7_u0_n171 ) , .A1( u2_u7_u0_n174 ) );
  NAND3_X1 u2_u7_u0_U93 (.A2( u2_u7_u0_n128 ) , .A1( u2_u7_u0_n132 ) , .A3( u2_u7_u0_n146 ) , .ZN( u2_u7_u0_n97 ) );
  OAI22_X1 u2_u7_u2_U10 (.ZN( u2_u7_u2_n109 ) , .A2( u2_u7_u2_n113 ) , .B2( u2_u7_u2_n133 ) , .B1( u2_u7_u2_n167 ) , .A1( u2_u7_u2_n168 ) );
  NAND3_X1 u2_u7_u2_U100 (.A2( u2_u7_u2_n100 ) , .A1( u2_u7_u2_n104 ) , .A3( u2_u7_u2_n138 ) , .ZN( u2_u7_u2_n98 ) );
  OAI22_X1 u2_u7_u2_U11 (.B1( u2_u7_u2_n151 ) , .A2( u2_u7_u2_n152 ) , .A1( u2_u7_u2_n153 ) , .ZN( u2_u7_u2_n160 ) , .B2( u2_u7_u2_n168 ) );
  NOR3_X1 u2_u7_u2_U12 (.A1( u2_u7_u2_n150 ) , .ZN( u2_u7_u2_n151 ) , .A3( u2_u7_u2_n175 ) , .A2( u2_u7_u2_n188 ) );
  AOI21_X1 u2_u7_u2_U13 (.ZN( u2_u7_u2_n144 ) , .B2( u2_u7_u2_n155 ) , .A( u2_u7_u2_n172 ) , .B1( u2_u7_u2_n185 ) );
  AOI21_X1 u2_u7_u2_U14 (.B2( u2_u7_u2_n143 ) , .ZN( u2_u7_u2_n145 ) , .B1( u2_u7_u2_n152 ) , .A( u2_u7_u2_n171 ) );
  AOI21_X1 u2_u7_u2_U15 (.B2( u2_u7_u2_n120 ) , .B1( u2_u7_u2_n121 ) , .ZN( u2_u7_u2_n126 ) , .A( u2_u7_u2_n167 ) );
  INV_X1 u2_u7_u2_U16 (.A( u2_u7_u2_n156 ) , .ZN( u2_u7_u2_n171 ) );
  INV_X1 u2_u7_u2_U17 (.A( u2_u7_u2_n120 ) , .ZN( u2_u7_u2_n188 ) );
  NAND2_X1 u2_u7_u2_U18 (.A2( u2_u7_u2_n122 ) , .ZN( u2_u7_u2_n150 ) , .A1( u2_u7_u2_n152 ) );
  INV_X1 u2_u7_u2_U19 (.A( u2_u7_u2_n153 ) , .ZN( u2_u7_u2_n170 ) );
  INV_X1 u2_u7_u2_U20 (.A( u2_u7_u2_n137 ) , .ZN( u2_u7_u2_n173 ) );
  NAND2_X1 u2_u7_u2_U21 (.A1( u2_u7_u2_n132 ) , .A2( u2_u7_u2_n139 ) , .ZN( u2_u7_u2_n157 ) );
  INV_X1 u2_u7_u2_U22 (.A( u2_u7_u2_n113 ) , .ZN( u2_u7_u2_n178 ) );
  INV_X1 u2_u7_u2_U23 (.A( u2_u7_u2_n139 ) , .ZN( u2_u7_u2_n175 ) );
  INV_X1 u2_u7_u2_U24 (.A( u2_u7_u2_n155 ) , .ZN( u2_u7_u2_n181 ) );
  INV_X1 u2_u7_u2_U25 (.A( u2_u7_u2_n119 ) , .ZN( u2_u7_u2_n177 ) );
  INV_X1 u2_u7_u2_U26 (.A( u2_u7_u2_n116 ) , .ZN( u2_u7_u2_n180 ) );
  INV_X1 u2_u7_u2_U27 (.A( u2_u7_u2_n131 ) , .ZN( u2_u7_u2_n179 ) );
  INV_X1 u2_u7_u2_U28 (.A( u2_u7_u2_n154 ) , .ZN( u2_u7_u2_n176 ) );
  NAND2_X1 u2_u7_u2_U29 (.A2( u2_u7_u2_n116 ) , .A1( u2_u7_u2_n117 ) , .ZN( u2_u7_u2_n118 ) );
  NOR2_X1 u2_u7_u2_U3 (.ZN( u2_u7_u2_n121 ) , .A2( u2_u7_u2_n177 ) , .A1( u2_u7_u2_n180 ) );
  INV_X1 u2_u7_u2_U30 (.A( u2_u7_u2_n132 ) , .ZN( u2_u7_u2_n182 ) );
  INV_X1 u2_u7_u2_U31 (.A( u2_u7_u2_n158 ) , .ZN( u2_u7_u2_n183 ) );
  OAI21_X1 u2_u7_u2_U32 (.A( u2_u7_u2_n156 ) , .B1( u2_u7_u2_n157 ) , .ZN( u2_u7_u2_n158 ) , .B2( u2_u7_u2_n179 ) );
  NOR2_X1 u2_u7_u2_U33 (.ZN( u2_u7_u2_n156 ) , .A1( u2_u7_u2_n166 ) , .A2( u2_u7_u2_n169 ) );
  NOR2_X1 u2_u7_u2_U34 (.A2( u2_u7_u2_n114 ) , .ZN( u2_u7_u2_n137 ) , .A1( u2_u7_u2_n140 ) );
  NOR2_X1 u2_u7_u2_U35 (.A2( u2_u7_u2_n138 ) , .ZN( u2_u7_u2_n153 ) , .A1( u2_u7_u2_n156 ) );
  AOI211_X1 u2_u7_u2_U36 (.ZN( u2_u7_u2_n130 ) , .C1( u2_u7_u2_n138 ) , .C2( u2_u7_u2_n179 ) , .B( u2_u7_u2_n96 ) , .A( u2_u7_u2_n97 ) );
  OAI22_X1 u2_u7_u2_U37 (.B1( u2_u7_u2_n133 ) , .A2( u2_u7_u2_n137 ) , .A1( u2_u7_u2_n152 ) , .B2( u2_u7_u2_n168 ) , .ZN( u2_u7_u2_n97 ) );
  OAI221_X1 u2_u7_u2_U38 (.B1( u2_u7_u2_n113 ) , .C1( u2_u7_u2_n132 ) , .A( u2_u7_u2_n149 ) , .B2( u2_u7_u2_n171 ) , .C2( u2_u7_u2_n172 ) , .ZN( u2_u7_u2_n96 ) );
  OAI221_X1 u2_u7_u2_U39 (.A( u2_u7_u2_n115 ) , .C2( u2_u7_u2_n123 ) , .B2( u2_u7_u2_n143 ) , .B1( u2_u7_u2_n153 ) , .ZN( u2_u7_u2_n163 ) , .C1( u2_u7_u2_n168 ) );
  INV_X1 u2_u7_u2_U4 (.A( u2_u7_u2_n134 ) , .ZN( u2_u7_u2_n185 ) );
  OAI21_X1 u2_u7_u2_U40 (.A( u2_u7_u2_n114 ) , .ZN( u2_u7_u2_n115 ) , .B1( u2_u7_u2_n176 ) , .B2( u2_u7_u2_n178 ) );
  OAI221_X1 u2_u7_u2_U41 (.A( u2_u7_u2_n135 ) , .B2( u2_u7_u2_n136 ) , .B1( u2_u7_u2_n137 ) , .ZN( u2_u7_u2_n162 ) , .C2( u2_u7_u2_n167 ) , .C1( u2_u7_u2_n185 ) );
  AND3_X1 u2_u7_u2_U42 (.A3( u2_u7_u2_n131 ) , .A2( u2_u7_u2_n132 ) , .A1( u2_u7_u2_n133 ) , .ZN( u2_u7_u2_n136 ) );
  AOI22_X1 u2_u7_u2_U43 (.ZN( u2_u7_u2_n135 ) , .B1( u2_u7_u2_n140 ) , .A1( u2_u7_u2_n156 ) , .B2( u2_u7_u2_n180 ) , .A2( u2_u7_u2_n188 ) );
  AOI21_X1 u2_u7_u2_U44 (.ZN( u2_u7_u2_n149 ) , .B1( u2_u7_u2_n173 ) , .B2( u2_u7_u2_n188 ) , .A( u2_u7_u2_n95 ) );
  AND3_X1 u2_u7_u2_U45 (.A2( u2_u7_u2_n100 ) , .A1( u2_u7_u2_n104 ) , .A3( u2_u7_u2_n156 ) , .ZN( u2_u7_u2_n95 ) );
  OAI21_X1 u2_u7_u2_U46 (.A( u2_u7_u2_n101 ) , .B2( u2_u7_u2_n121 ) , .B1( u2_u7_u2_n153 ) , .ZN( u2_u7_u2_n164 ) );
  NAND2_X1 u2_u7_u2_U47 (.A2( u2_u7_u2_n100 ) , .A1( u2_u7_u2_n107 ) , .ZN( u2_u7_u2_n155 ) );
  NAND2_X1 u2_u7_u2_U48 (.A2( u2_u7_u2_n105 ) , .A1( u2_u7_u2_n108 ) , .ZN( u2_u7_u2_n143 ) );
  NAND2_X1 u2_u7_u2_U49 (.A1( u2_u7_u2_n104 ) , .A2( u2_u7_u2_n106 ) , .ZN( u2_u7_u2_n152 ) );
  INV_X1 u2_u7_u2_U5 (.A( u2_u7_u2_n150 ) , .ZN( u2_u7_u2_n184 ) );
  NAND2_X1 u2_u7_u2_U50 (.A1( u2_u7_u2_n100 ) , .A2( u2_u7_u2_n105 ) , .ZN( u2_u7_u2_n132 ) );
  INV_X1 u2_u7_u2_U51 (.A( u2_u7_u2_n140 ) , .ZN( u2_u7_u2_n168 ) );
  INV_X1 u2_u7_u2_U52 (.A( u2_u7_u2_n138 ) , .ZN( u2_u7_u2_n167 ) );
  OAI21_X1 u2_u7_u2_U53 (.A( u2_u7_u2_n141 ) , .B2( u2_u7_u2_n142 ) , .ZN( u2_u7_u2_n146 ) , .B1( u2_u7_u2_n153 ) );
  OAI21_X1 u2_u7_u2_U54 (.A( u2_u7_u2_n140 ) , .ZN( u2_u7_u2_n141 ) , .B1( u2_u7_u2_n176 ) , .B2( u2_u7_u2_n177 ) );
  NOR3_X1 u2_u7_u2_U55 (.ZN( u2_u7_u2_n142 ) , .A3( u2_u7_u2_n175 ) , .A2( u2_u7_u2_n178 ) , .A1( u2_u7_u2_n181 ) );
  INV_X1 u2_u7_u2_U56 (.ZN( u2_u7_u2_n187 ) , .A( u2_u7_u2_n99 ) );
  OAI21_X1 u2_u7_u2_U57 (.B1( u2_u7_u2_n137 ) , .B2( u2_u7_u2_n143 ) , .A( u2_u7_u2_n98 ) , .ZN( u2_u7_u2_n99 ) );
  NAND2_X1 u2_u7_u2_U58 (.A1( u2_u7_u2_n102 ) , .A2( u2_u7_u2_n106 ) , .ZN( u2_u7_u2_n113 ) );
  NAND2_X1 u2_u7_u2_U59 (.A1( u2_u7_u2_n106 ) , .A2( u2_u7_u2_n107 ) , .ZN( u2_u7_u2_n131 ) );
  NOR4_X1 u2_u7_u2_U6 (.A4( u2_u7_u2_n124 ) , .A3( u2_u7_u2_n125 ) , .A2( u2_u7_u2_n126 ) , .A1( u2_u7_u2_n127 ) , .ZN( u2_u7_u2_n128 ) );
  NAND2_X1 u2_u7_u2_U60 (.A1( u2_u7_u2_n103 ) , .A2( u2_u7_u2_n107 ) , .ZN( u2_u7_u2_n139 ) );
  NAND2_X1 u2_u7_u2_U61 (.A1( u2_u7_u2_n103 ) , .A2( u2_u7_u2_n105 ) , .ZN( u2_u7_u2_n133 ) );
  NAND2_X1 u2_u7_u2_U62 (.A1( u2_u7_u2_n102 ) , .A2( u2_u7_u2_n103 ) , .ZN( u2_u7_u2_n154 ) );
  NAND2_X1 u2_u7_u2_U63 (.A2( u2_u7_u2_n103 ) , .A1( u2_u7_u2_n104 ) , .ZN( u2_u7_u2_n119 ) );
  NAND2_X1 u2_u7_u2_U64 (.A2( u2_u7_u2_n107 ) , .A1( u2_u7_u2_n108 ) , .ZN( u2_u7_u2_n123 ) );
  NAND2_X1 u2_u7_u2_U65 (.A1( u2_u7_u2_n104 ) , .A2( u2_u7_u2_n108 ) , .ZN( u2_u7_u2_n122 ) );
  INV_X1 u2_u7_u2_U66 (.A( u2_u7_u2_n114 ) , .ZN( u2_u7_u2_n172 ) );
  NAND2_X1 u2_u7_u2_U67 (.A2( u2_u7_u2_n100 ) , .A1( u2_u7_u2_n102 ) , .ZN( u2_u7_u2_n116 ) );
  NAND2_X1 u2_u7_u2_U68 (.A1( u2_u7_u2_n102 ) , .A2( u2_u7_u2_n108 ) , .ZN( u2_u7_u2_n120 ) );
  NAND2_X1 u2_u7_u2_U69 (.A2( u2_u7_u2_n105 ) , .A1( u2_u7_u2_n106 ) , .ZN( u2_u7_u2_n117 ) );
  AOI21_X1 u2_u7_u2_U7 (.B2( u2_u7_u2_n119 ) , .ZN( u2_u7_u2_n127 ) , .A( u2_u7_u2_n137 ) , .B1( u2_u7_u2_n155 ) );
  NOR2_X1 u2_u7_u2_U70 (.A2( u2_u7_X_16 ) , .ZN( u2_u7_u2_n140 ) , .A1( u2_u7_u2_n166 ) );
  NOR2_X1 u2_u7_u2_U71 (.A2( u2_u7_X_13 ) , .A1( u2_u7_X_14 ) , .ZN( u2_u7_u2_n100 ) );
  NOR2_X1 u2_u7_u2_U72 (.A2( u2_u7_X_16 ) , .A1( u2_u7_X_17 ) , .ZN( u2_u7_u2_n138 ) );
  NOR2_X1 u2_u7_u2_U73 (.A2( u2_u7_X_15 ) , .A1( u2_u7_X_18 ) , .ZN( u2_u7_u2_n104 ) );
  NOR2_X1 u2_u7_u2_U74 (.A2( u2_u7_X_14 ) , .ZN( u2_u7_u2_n103 ) , .A1( u2_u7_u2_n174 ) );
  NOR2_X1 u2_u7_u2_U75 (.A2( u2_u7_X_15 ) , .ZN( u2_u7_u2_n102 ) , .A1( u2_u7_u2_n165 ) );
  NOR2_X1 u2_u7_u2_U76 (.A2( u2_u7_X_17 ) , .ZN( u2_u7_u2_n114 ) , .A1( u2_u7_u2_n169 ) );
  AND2_X1 u2_u7_u2_U77 (.A1( u2_u7_X_15 ) , .ZN( u2_u7_u2_n105 ) , .A2( u2_u7_u2_n165 ) );
  AND2_X1 u2_u7_u2_U78 (.A2( u2_u7_X_15 ) , .A1( u2_u7_X_18 ) , .ZN( u2_u7_u2_n107 ) );
  AND2_X1 u2_u7_u2_U79 (.A1( u2_u7_X_14 ) , .ZN( u2_u7_u2_n106 ) , .A2( u2_u7_u2_n174 ) );
  AOI21_X1 u2_u7_u2_U8 (.ZN( u2_u7_u2_n124 ) , .B1( u2_u7_u2_n131 ) , .B2( u2_u7_u2_n143 ) , .A( u2_u7_u2_n172 ) );
  AND2_X1 u2_u7_u2_U80 (.A1( u2_u7_X_13 ) , .A2( u2_u7_X_14 ) , .ZN( u2_u7_u2_n108 ) );
  INV_X1 u2_u7_u2_U81 (.A( u2_u7_X_16 ) , .ZN( u2_u7_u2_n169 ) );
  INV_X1 u2_u7_u2_U82 (.A( u2_u7_X_17 ) , .ZN( u2_u7_u2_n166 ) );
  INV_X1 u2_u7_u2_U83 (.A( u2_u7_X_13 ) , .ZN( u2_u7_u2_n174 ) );
  INV_X1 u2_u7_u2_U84 (.A( u2_u7_X_18 ) , .ZN( u2_u7_u2_n165 ) );
  NAND4_X1 u2_u7_u2_U85 (.ZN( u2_out7_24 ) , .A4( u2_u7_u2_n111 ) , .A3( u2_u7_u2_n112 ) , .A1( u2_u7_u2_n130 ) , .A2( u2_u7_u2_n187 ) );
  AOI221_X1 u2_u7_u2_U86 (.A( u2_u7_u2_n109 ) , .B1( u2_u7_u2_n110 ) , .ZN( u2_u7_u2_n111 ) , .C1( u2_u7_u2_n134 ) , .C2( u2_u7_u2_n170 ) , .B2( u2_u7_u2_n173 ) );
  AOI21_X1 u2_u7_u2_U87 (.ZN( u2_u7_u2_n112 ) , .B2( u2_u7_u2_n156 ) , .A( u2_u7_u2_n164 ) , .B1( u2_u7_u2_n181 ) );
  NAND4_X1 u2_u7_u2_U88 (.ZN( u2_out7_16 ) , .A4( u2_u7_u2_n128 ) , .A3( u2_u7_u2_n129 ) , .A1( u2_u7_u2_n130 ) , .A2( u2_u7_u2_n186 ) );
  AOI22_X1 u2_u7_u2_U89 (.A2( u2_u7_u2_n118 ) , .ZN( u2_u7_u2_n129 ) , .A1( u2_u7_u2_n140 ) , .B1( u2_u7_u2_n157 ) , .B2( u2_u7_u2_n170 ) );
  AOI21_X1 u2_u7_u2_U9 (.B2( u2_u7_u2_n123 ) , .ZN( u2_u7_u2_n125 ) , .A( u2_u7_u2_n171 ) , .B1( u2_u7_u2_n184 ) );
  INV_X1 u2_u7_u2_U90 (.A( u2_u7_u2_n163 ) , .ZN( u2_u7_u2_n186 ) );
  NAND4_X1 u2_u7_u2_U91 (.ZN( u2_out7_30 ) , .A4( u2_u7_u2_n147 ) , .A3( u2_u7_u2_n148 ) , .A2( u2_u7_u2_n149 ) , .A1( u2_u7_u2_n187 ) );
  NOR3_X1 u2_u7_u2_U92 (.A3( u2_u7_u2_n144 ) , .A2( u2_u7_u2_n145 ) , .A1( u2_u7_u2_n146 ) , .ZN( u2_u7_u2_n147 ) );
  AOI21_X1 u2_u7_u2_U93 (.B2( u2_u7_u2_n138 ) , .ZN( u2_u7_u2_n148 ) , .A( u2_u7_u2_n162 ) , .B1( u2_u7_u2_n182 ) );
  OR4_X1 u2_u7_u2_U94 (.ZN( u2_out7_6 ) , .A4( u2_u7_u2_n161 ) , .A3( u2_u7_u2_n162 ) , .A2( u2_u7_u2_n163 ) , .A1( u2_u7_u2_n164 ) );
  OR3_X1 u2_u7_u2_U95 (.A2( u2_u7_u2_n159 ) , .A1( u2_u7_u2_n160 ) , .ZN( u2_u7_u2_n161 ) , .A3( u2_u7_u2_n183 ) );
  AOI21_X1 u2_u7_u2_U96 (.B2( u2_u7_u2_n154 ) , .B1( u2_u7_u2_n155 ) , .ZN( u2_u7_u2_n159 ) , .A( u2_u7_u2_n167 ) );
  NAND3_X1 u2_u7_u2_U97 (.A2( u2_u7_u2_n117 ) , .A1( u2_u7_u2_n122 ) , .A3( u2_u7_u2_n123 ) , .ZN( u2_u7_u2_n134 ) );
  NAND3_X1 u2_u7_u2_U98 (.ZN( u2_u7_u2_n110 ) , .A2( u2_u7_u2_n131 ) , .A3( u2_u7_u2_n139 ) , .A1( u2_u7_u2_n154 ) );
  NAND3_X1 u2_u7_u2_U99 (.A2( u2_u7_u2_n100 ) , .ZN( u2_u7_u2_n101 ) , .A1( u2_u7_u2_n104 ) , .A3( u2_u7_u2_n114 ) );
  XOR2_X1 u2_u8_U26 (.B( u2_K9_30 ) , .A( u2_R7_21 ) , .Z( u2_u8_X_30 ) );
  XOR2_X1 u2_u8_U28 (.B( u2_K9_29 ) , .A( u2_R7_20 ) , .Z( u2_u8_X_29 ) );
  XOR2_X1 u2_u8_U29 (.B( u2_K9_28 ) , .A( u2_R7_19 ) , .Z( u2_u8_X_28 ) );
  XOR2_X1 u2_u8_U30 (.B( u2_K9_27 ) , .A( u2_R7_18 ) , .Z( u2_u8_X_27 ) );
  XOR2_X1 u2_u8_U31 (.B( u2_K9_26 ) , .A( u2_R7_17 ) , .Z( u2_u8_X_26 ) );
  XOR2_X1 u2_u8_U32 (.B( u2_K9_25 ) , .A( u2_R7_16 ) , .Z( u2_u8_X_25 ) );
  XOR2_X1 u2_u8_U33 (.B( u2_K9_24 ) , .A( u2_R7_17 ) , .Z( u2_u8_X_24 ) );
  XOR2_X1 u2_u8_U34 (.B( u2_K9_23 ) , .A( u2_R7_16 ) , .Z( u2_u8_X_23 ) );
  XOR2_X1 u2_u8_U35 (.B( u2_K9_22 ) , .A( u2_R7_15 ) , .Z( u2_u8_X_22 ) );
  XOR2_X1 u2_u8_U36 (.B( u2_K9_21 ) , .A( u2_R7_14 ) , .Z( u2_u8_X_21 ) );
  XOR2_X1 u2_u8_U37 (.B( u2_K9_20 ) , .A( u2_R7_13 ) , .Z( u2_u8_X_20 ) );
  XOR2_X1 u2_u8_U39 (.B( u2_K9_19 ) , .A( u2_R7_12 ) , .Z( u2_u8_X_19 ) );
  OAI22_X1 u2_u8_u3_U10 (.B1( u2_u8_u3_n113 ) , .A2( u2_u8_u3_n135 ) , .A1( u2_u8_u3_n150 ) , .B2( u2_u8_u3_n164 ) , .ZN( u2_u8_u3_n98 ) );
  OAI211_X1 u2_u8_u3_U11 (.B( u2_u8_u3_n106 ) , .ZN( u2_u8_u3_n119 ) , .C2( u2_u8_u3_n128 ) , .C1( u2_u8_u3_n167 ) , .A( u2_u8_u3_n181 ) );
  AOI221_X1 u2_u8_u3_U12 (.C1( u2_u8_u3_n105 ) , .ZN( u2_u8_u3_n106 ) , .A( u2_u8_u3_n131 ) , .B2( u2_u8_u3_n132 ) , .C2( u2_u8_u3_n133 ) , .B1( u2_u8_u3_n169 ) );
  INV_X1 u2_u8_u3_U13 (.ZN( u2_u8_u3_n181 ) , .A( u2_u8_u3_n98 ) );
  NAND2_X1 u2_u8_u3_U14 (.ZN( u2_u8_u3_n105 ) , .A2( u2_u8_u3_n130 ) , .A1( u2_u8_u3_n155 ) );
  AOI22_X1 u2_u8_u3_U15 (.B1( u2_u8_u3_n115 ) , .A2( u2_u8_u3_n116 ) , .ZN( u2_u8_u3_n123 ) , .B2( u2_u8_u3_n133 ) , .A1( u2_u8_u3_n169 ) );
  NAND2_X1 u2_u8_u3_U16 (.ZN( u2_u8_u3_n116 ) , .A2( u2_u8_u3_n151 ) , .A1( u2_u8_u3_n182 ) );
  NOR2_X1 u2_u8_u3_U17 (.ZN( u2_u8_u3_n126 ) , .A2( u2_u8_u3_n150 ) , .A1( u2_u8_u3_n164 ) );
  AOI21_X1 u2_u8_u3_U18 (.ZN( u2_u8_u3_n112 ) , .B2( u2_u8_u3_n146 ) , .B1( u2_u8_u3_n155 ) , .A( u2_u8_u3_n167 ) );
  NAND2_X1 u2_u8_u3_U19 (.A1( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n142 ) , .A2( u2_u8_u3_n164 ) );
  NAND2_X1 u2_u8_u3_U20 (.ZN( u2_u8_u3_n132 ) , .A2( u2_u8_u3_n152 ) , .A1( u2_u8_u3_n156 ) );
  AND2_X1 u2_u8_u3_U21 (.A2( u2_u8_u3_n113 ) , .A1( u2_u8_u3_n114 ) , .ZN( u2_u8_u3_n151 ) );
  INV_X1 u2_u8_u3_U22 (.A( u2_u8_u3_n133 ) , .ZN( u2_u8_u3_n165 ) );
  INV_X1 u2_u8_u3_U23 (.A( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n170 ) );
  NAND2_X1 u2_u8_u3_U24 (.A1( u2_u8_u3_n107 ) , .A2( u2_u8_u3_n108 ) , .ZN( u2_u8_u3_n140 ) );
  NAND2_X1 u2_u8_u3_U25 (.ZN( u2_u8_u3_n117 ) , .A1( u2_u8_u3_n124 ) , .A2( u2_u8_u3_n148 ) );
  NAND2_X1 u2_u8_u3_U26 (.ZN( u2_u8_u3_n143 ) , .A1( u2_u8_u3_n165 ) , .A2( u2_u8_u3_n167 ) );
  INV_X1 u2_u8_u3_U27 (.A( u2_u8_u3_n130 ) , .ZN( u2_u8_u3_n177 ) );
  INV_X1 u2_u8_u3_U28 (.A( u2_u8_u3_n128 ) , .ZN( u2_u8_u3_n176 ) );
  INV_X1 u2_u8_u3_U29 (.A( u2_u8_u3_n155 ) , .ZN( u2_u8_u3_n174 ) );
  INV_X1 u2_u8_u3_U3 (.A( u2_u8_u3_n129 ) , .ZN( u2_u8_u3_n183 ) );
  INV_X1 u2_u8_u3_U30 (.A( u2_u8_u3_n139 ) , .ZN( u2_u8_u3_n185 ) );
  NOR2_X1 u2_u8_u3_U31 (.ZN( u2_u8_u3_n135 ) , .A2( u2_u8_u3_n141 ) , .A1( u2_u8_u3_n169 ) );
  OAI222_X1 u2_u8_u3_U32 (.C2( u2_u8_u3_n107 ) , .A2( u2_u8_u3_n108 ) , .B1( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n138 ) , .B2( u2_u8_u3_n146 ) , .C1( u2_u8_u3_n154 ) , .A1( u2_u8_u3_n164 ) );
  NOR4_X1 u2_u8_u3_U33 (.A4( u2_u8_u3_n157 ) , .A3( u2_u8_u3_n158 ) , .A2( u2_u8_u3_n159 ) , .A1( u2_u8_u3_n160 ) , .ZN( u2_u8_u3_n161 ) );
  AOI21_X1 u2_u8_u3_U34 (.B2( u2_u8_u3_n152 ) , .B1( u2_u8_u3_n153 ) , .ZN( u2_u8_u3_n158 ) , .A( u2_u8_u3_n164 ) );
  AOI21_X1 u2_u8_u3_U35 (.A( u2_u8_u3_n149 ) , .B2( u2_u8_u3_n150 ) , .B1( u2_u8_u3_n151 ) , .ZN( u2_u8_u3_n159 ) );
  AOI21_X1 u2_u8_u3_U36 (.A( u2_u8_u3_n154 ) , .B2( u2_u8_u3_n155 ) , .B1( u2_u8_u3_n156 ) , .ZN( u2_u8_u3_n157 ) );
  AOI211_X1 u2_u8_u3_U37 (.ZN( u2_u8_u3_n109 ) , .A( u2_u8_u3_n119 ) , .C2( u2_u8_u3_n129 ) , .B( u2_u8_u3_n138 ) , .C1( u2_u8_u3_n141 ) );
  AOI211_X1 u2_u8_u3_U38 (.B( u2_u8_u3_n119 ) , .A( u2_u8_u3_n120 ) , .C2( u2_u8_u3_n121 ) , .ZN( u2_u8_u3_n122 ) , .C1( u2_u8_u3_n179 ) );
  INV_X1 u2_u8_u3_U39 (.A( u2_u8_u3_n156 ) , .ZN( u2_u8_u3_n179 ) );
  INV_X1 u2_u8_u3_U4 (.A( u2_u8_u3_n140 ) , .ZN( u2_u8_u3_n182 ) );
  OAI22_X1 u2_u8_u3_U40 (.B1( u2_u8_u3_n118 ) , .ZN( u2_u8_u3_n120 ) , .A1( u2_u8_u3_n135 ) , .B2( u2_u8_u3_n154 ) , .A2( u2_u8_u3_n178 ) );
  AND3_X1 u2_u8_u3_U41 (.ZN( u2_u8_u3_n118 ) , .A2( u2_u8_u3_n124 ) , .A1( u2_u8_u3_n144 ) , .A3( u2_u8_u3_n152 ) );
  INV_X1 u2_u8_u3_U42 (.A( u2_u8_u3_n121 ) , .ZN( u2_u8_u3_n164 ) );
  NAND2_X1 u2_u8_u3_U43 (.ZN( u2_u8_u3_n133 ) , .A1( u2_u8_u3_n154 ) , .A2( u2_u8_u3_n164 ) );
  OAI211_X1 u2_u8_u3_U44 (.B( u2_u8_u3_n127 ) , .ZN( u2_u8_u3_n139 ) , .C1( u2_u8_u3_n150 ) , .C2( u2_u8_u3_n154 ) , .A( u2_u8_u3_n184 ) );
  INV_X1 u2_u8_u3_U45 (.A( u2_u8_u3_n125 ) , .ZN( u2_u8_u3_n184 ) );
  AOI221_X1 u2_u8_u3_U46 (.A( u2_u8_u3_n126 ) , .ZN( u2_u8_u3_n127 ) , .C2( u2_u8_u3_n132 ) , .C1( u2_u8_u3_n169 ) , .B2( u2_u8_u3_n170 ) , .B1( u2_u8_u3_n174 ) );
  OAI22_X1 u2_u8_u3_U47 (.A1( u2_u8_u3_n124 ) , .ZN( u2_u8_u3_n125 ) , .B2( u2_u8_u3_n145 ) , .A2( u2_u8_u3_n165 ) , .B1( u2_u8_u3_n167 ) );
  NOR2_X1 u2_u8_u3_U48 (.A1( u2_u8_u3_n113 ) , .ZN( u2_u8_u3_n131 ) , .A2( u2_u8_u3_n154 ) );
  NAND2_X1 u2_u8_u3_U49 (.A1( u2_u8_u3_n103 ) , .ZN( u2_u8_u3_n150 ) , .A2( u2_u8_u3_n99 ) );
  INV_X1 u2_u8_u3_U5 (.A( u2_u8_u3_n117 ) , .ZN( u2_u8_u3_n178 ) );
  NAND2_X1 u2_u8_u3_U50 (.A2( u2_u8_u3_n102 ) , .ZN( u2_u8_u3_n155 ) , .A1( u2_u8_u3_n97 ) );
  INV_X1 u2_u8_u3_U51 (.A( u2_u8_u3_n141 ) , .ZN( u2_u8_u3_n167 ) );
  AOI21_X1 u2_u8_u3_U52 (.B2( u2_u8_u3_n114 ) , .B1( u2_u8_u3_n146 ) , .A( u2_u8_u3_n154 ) , .ZN( u2_u8_u3_n94 ) );
  AOI21_X1 u2_u8_u3_U53 (.ZN( u2_u8_u3_n110 ) , .B2( u2_u8_u3_n142 ) , .B1( u2_u8_u3_n186 ) , .A( u2_u8_u3_n95 ) );
  INV_X1 u2_u8_u3_U54 (.A( u2_u8_u3_n145 ) , .ZN( u2_u8_u3_n186 ) );
  AOI21_X1 u2_u8_u3_U55 (.B1( u2_u8_u3_n124 ) , .A( u2_u8_u3_n149 ) , .B2( u2_u8_u3_n155 ) , .ZN( u2_u8_u3_n95 ) );
  INV_X1 u2_u8_u3_U56 (.A( u2_u8_u3_n149 ) , .ZN( u2_u8_u3_n169 ) );
  NAND2_X1 u2_u8_u3_U57 (.ZN( u2_u8_u3_n124 ) , .A1( u2_u8_u3_n96 ) , .A2( u2_u8_u3_n97 ) );
  NAND2_X1 u2_u8_u3_U58 (.A2( u2_u8_u3_n100 ) , .ZN( u2_u8_u3_n146 ) , .A1( u2_u8_u3_n96 ) );
  NAND2_X1 u2_u8_u3_U59 (.A1( u2_u8_u3_n101 ) , .ZN( u2_u8_u3_n145 ) , .A2( u2_u8_u3_n99 ) );
  AOI221_X1 u2_u8_u3_U6 (.A( u2_u8_u3_n131 ) , .C2( u2_u8_u3_n132 ) , .C1( u2_u8_u3_n133 ) , .ZN( u2_u8_u3_n134 ) , .B1( u2_u8_u3_n143 ) , .B2( u2_u8_u3_n177 ) );
  NAND2_X1 u2_u8_u3_U60 (.A1( u2_u8_u3_n100 ) , .ZN( u2_u8_u3_n156 ) , .A2( u2_u8_u3_n99 ) );
  NAND2_X1 u2_u8_u3_U61 (.A2( u2_u8_u3_n101 ) , .A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n148 ) );
  NAND2_X1 u2_u8_u3_U62 (.A1( u2_u8_u3_n100 ) , .A2( u2_u8_u3_n102 ) , .ZN( u2_u8_u3_n128 ) );
  NAND2_X1 u2_u8_u3_U63 (.A2( u2_u8_u3_n101 ) , .A1( u2_u8_u3_n102 ) , .ZN( u2_u8_u3_n152 ) );
  NAND2_X1 u2_u8_u3_U64 (.A2( u2_u8_u3_n101 ) , .ZN( u2_u8_u3_n114 ) , .A1( u2_u8_u3_n96 ) );
  NAND2_X1 u2_u8_u3_U65 (.ZN( u2_u8_u3_n107 ) , .A1( u2_u8_u3_n97 ) , .A2( u2_u8_u3_n99 ) );
  NAND2_X1 u2_u8_u3_U66 (.A2( u2_u8_u3_n100 ) , .A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n113 ) );
  NAND2_X1 u2_u8_u3_U67 (.A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n153 ) , .A2( u2_u8_u3_n97 ) );
  NAND2_X1 u2_u8_u3_U68 (.A2( u2_u8_u3_n103 ) , .A1( u2_u8_u3_n104 ) , .ZN( u2_u8_u3_n130 ) );
  NAND2_X1 u2_u8_u3_U69 (.A2( u2_u8_u3_n103 ) , .ZN( u2_u8_u3_n144 ) , .A1( u2_u8_u3_n96 ) );
  OAI22_X1 u2_u8_u3_U7 (.B2( u2_u8_u3_n147 ) , .A2( u2_u8_u3_n148 ) , .ZN( u2_u8_u3_n160 ) , .B1( u2_u8_u3_n165 ) , .A1( u2_u8_u3_n168 ) );
  NAND2_X1 u2_u8_u3_U70 (.A1( u2_u8_u3_n102 ) , .A2( u2_u8_u3_n103 ) , .ZN( u2_u8_u3_n108 ) );
  NOR2_X1 u2_u8_u3_U71 (.A2( u2_u8_X_19 ) , .A1( u2_u8_X_20 ) , .ZN( u2_u8_u3_n99 ) );
  NOR2_X1 u2_u8_u3_U72 (.A2( u2_u8_X_21 ) , .A1( u2_u8_X_24 ) , .ZN( u2_u8_u3_n103 ) );
  NOR2_X1 u2_u8_u3_U73 (.A2( u2_u8_X_24 ) , .A1( u2_u8_u3_n171 ) , .ZN( u2_u8_u3_n97 ) );
  NOR2_X1 u2_u8_u3_U74 (.A2( u2_u8_X_23 ) , .ZN( u2_u8_u3_n141 ) , .A1( u2_u8_u3_n166 ) );
  NOR2_X1 u2_u8_u3_U75 (.A2( u2_u8_X_19 ) , .A1( u2_u8_u3_n172 ) , .ZN( u2_u8_u3_n96 ) );
  NAND2_X1 u2_u8_u3_U76 (.A1( u2_u8_X_22 ) , .A2( u2_u8_X_23 ) , .ZN( u2_u8_u3_n154 ) );
  NAND2_X1 u2_u8_u3_U77 (.A1( u2_u8_X_23 ) , .ZN( u2_u8_u3_n149 ) , .A2( u2_u8_u3_n166 ) );
  NOR2_X1 u2_u8_u3_U78 (.A2( u2_u8_X_22 ) , .A1( u2_u8_X_23 ) , .ZN( u2_u8_u3_n121 ) );
  AND2_X1 u2_u8_u3_U79 (.A1( u2_u8_X_24 ) , .ZN( u2_u8_u3_n101 ) , .A2( u2_u8_u3_n171 ) );
  AND3_X1 u2_u8_u3_U8 (.A3( u2_u8_u3_n144 ) , .A2( u2_u8_u3_n145 ) , .A1( u2_u8_u3_n146 ) , .ZN( u2_u8_u3_n147 ) );
  AND2_X1 u2_u8_u3_U80 (.A1( u2_u8_X_19 ) , .ZN( u2_u8_u3_n102 ) , .A2( u2_u8_u3_n172 ) );
  AND2_X1 u2_u8_u3_U81 (.A1( u2_u8_X_21 ) , .A2( u2_u8_X_24 ) , .ZN( u2_u8_u3_n100 ) );
  AND2_X1 u2_u8_u3_U82 (.A2( u2_u8_X_19 ) , .A1( u2_u8_X_20 ) , .ZN( u2_u8_u3_n104 ) );
  INV_X1 u2_u8_u3_U83 (.A( u2_u8_X_22 ) , .ZN( u2_u8_u3_n166 ) );
  INV_X1 u2_u8_u3_U84 (.A( u2_u8_X_21 ) , .ZN( u2_u8_u3_n171 ) );
  INV_X1 u2_u8_u3_U85 (.A( u2_u8_X_20 ) , .ZN( u2_u8_u3_n172 ) );
  OR4_X1 u2_u8_u3_U86 (.ZN( u2_out8_10 ) , .A4( u2_u8_u3_n136 ) , .A3( u2_u8_u3_n137 ) , .A1( u2_u8_u3_n138 ) , .A2( u2_u8_u3_n139 ) );
  OAI222_X1 u2_u8_u3_U87 (.C1( u2_u8_u3_n128 ) , .ZN( u2_u8_u3_n137 ) , .B1( u2_u8_u3_n148 ) , .A2( u2_u8_u3_n150 ) , .B2( u2_u8_u3_n154 ) , .C2( u2_u8_u3_n164 ) , .A1( u2_u8_u3_n167 ) );
  OAI221_X1 u2_u8_u3_U88 (.A( u2_u8_u3_n134 ) , .B2( u2_u8_u3_n135 ) , .ZN( u2_u8_u3_n136 ) , .C1( u2_u8_u3_n149 ) , .B1( u2_u8_u3_n151 ) , .C2( u2_u8_u3_n183 ) );
  NAND4_X1 u2_u8_u3_U89 (.ZN( u2_out8_26 ) , .A4( u2_u8_u3_n109 ) , .A3( u2_u8_u3_n110 ) , .A2( u2_u8_u3_n111 ) , .A1( u2_u8_u3_n173 ) );
  INV_X1 u2_u8_u3_U9 (.A( u2_u8_u3_n143 ) , .ZN( u2_u8_u3_n168 ) );
  INV_X1 u2_u8_u3_U90 (.ZN( u2_u8_u3_n173 ) , .A( u2_u8_u3_n94 ) );
  OAI21_X1 u2_u8_u3_U91 (.ZN( u2_u8_u3_n111 ) , .B2( u2_u8_u3_n117 ) , .A( u2_u8_u3_n133 ) , .B1( u2_u8_u3_n176 ) );
  NAND4_X1 u2_u8_u3_U92 (.ZN( u2_out8_20 ) , .A4( u2_u8_u3_n122 ) , .A3( u2_u8_u3_n123 ) , .A1( u2_u8_u3_n175 ) , .A2( u2_u8_u3_n180 ) );
  INV_X1 u2_u8_u3_U93 (.A( u2_u8_u3_n126 ) , .ZN( u2_u8_u3_n180 ) );
  INV_X1 u2_u8_u3_U94 (.A( u2_u8_u3_n112 ) , .ZN( u2_u8_u3_n175 ) );
  NAND4_X1 u2_u8_u3_U95 (.ZN( u2_out8_1 ) , .A4( u2_u8_u3_n161 ) , .A3( u2_u8_u3_n162 ) , .A2( u2_u8_u3_n163 ) , .A1( u2_u8_u3_n185 ) );
  NAND2_X1 u2_u8_u3_U96 (.ZN( u2_u8_u3_n163 ) , .A2( u2_u8_u3_n170 ) , .A1( u2_u8_u3_n176 ) );
  AOI22_X1 u2_u8_u3_U97 (.B2( u2_u8_u3_n140 ) , .B1( u2_u8_u3_n141 ) , .A2( u2_u8_u3_n142 ) , .ZN( u2_u8_u3_n162 ) , .A1( u2_u8_u3_n177 ) );
  NAND3_X1 u2_u8_u3_U98 (.A1( u2_u8_u3_n114 ) , .ZN( u2_u8_u3_n115 ) , .A2( u2_u8_u3_n145 ) , .A3( u2_u8_u3_n153 ) );
  NAND3_X1 u2_u8_u3_U99 (.ZN( u2_u8_u3_n129 ) , .A2( u2_u8_u3_n144 ) , .A1( u2_u8_u3_n153 ) , .A3( u2_u8_u3_n182 ) );
  OAI22_X1 u2_u8_u4_U10 (.B2( u2_u8_u4_n135 ) , .ZN( u2_u8_u4_n137 ) , .B1( u2_u8_u4_n153 ) , .A1( u2_u8_u4_n155 ) , .A2( u2_u8_u4_n171 ) );
  AND3_X1 u2_u8_u4_U11 (.A2( u2_u8_u4_n134 ) , .ZN( u2_u8_u4_n135 ) , .A3( u2_u8_u4_n145 ) , .A1( u2_u8_u4_n157 ) );
  NAND2_X1 u2_u8_u4_U12 (.ZN( u2_u8_u4_n132 ) , .A2( u2_u8_u4_n170 ) , .A1( u2_u8_u4_n173 ) );
  AOI21_X1 u2_u8_u4_U13 (.B2( u2_u8_u4_n160 ) , .B1( u2_u8_u4_n161 ) , .ZN( u2_u8_u4_n162 ) , .A( u2_u8_u4_n170 ) );
  AOI21_X1 u2_u8_u4_U14 (.ZN( u2_u8_u4_n107 ) , .B2( u2_u8_u4_n143 ) , .A( u2_u8_u4_n174 ) , .B1( u2_u8_u4_n184 ) );
  AOI21_X1 u2_u8_u4_U15 (.B2( u2_u8_u4_n158 ) , .B1( u2_u8_u4_n159 ) , .ZN( u2_u8_u4_n163 ) , .A( u2_u8_u4_n174 ) );
  AOI21_X1 u2_u8_u4_U16 (.A( u2_u8_u4_n153 ) , .B2( u2_u8_u4_n154 ) , .B1( u2_u8_u4_n155 ) , .ZN( u2_u8_u4_n165 ) );
  AOI21_X1 u2_u8_u4_U17 (.A( u2_u8_u4_n156 ) , .B2( u2_u8_u4_n157 ) , .ZN( u2_u8_u4_n164 ) , .B1( u2_u8_u4_n184 ) );
  INV_X1 u2_u8_u4_U18 (.A( u2_u8_u4_n138 ) , .ZN( u2_u8_u4_n170 ) );
  AND2_X1 u2_u8_u4_U19 (.A2( u2_u8_u4_n120 ) , .ZN( u2_u8_u4_n155 ) , .A1( u2_u8_u4_n160 ) );
  INV_X1 u2_u8_u4_U20 (.A( u2_u8_u4_n156 ) , .ZN( u2_u8_u4_n175 ) );
  NAND2_X1 u2_u8_u4_U21 (.A2( u2_u8_u4_n118 ) , .ZN( u2_u8_u4_n131 ) , .A1( u2_u8_u4_n147 ) );
  NAND2_X1 u2_u8_u4_U22 (.A1( u2_u8_u4_n119 ) , .A2( u2_u8_u4_n120 ) , .ZN( u2_u8_u4_n130 ) );
  NAND2_X1 u2_u8_u4_U23 (.ZN( u2_u8_u4_n117 ) , .A2( u2_u8_u4_n118 ) , .A1( u2_u8_u4_n148 ) );
  NAND2_X1 u2_u8_u4_U24 (.ZN( u2_u8_u4_n129 ) , .A1( u2_u8_u4_n134 ) , .A2( u2_u8_u4_n148 ) );
  AND3_X1 u2_u8_u4_U25 (.A1( u2_u8_u4_n119 ) , .A2( u2_u8_u4_n143 ) , .A3( u2_u8_u4_n154 ) , .ZN( u2_u8_u4_n161 ) );
  AND2_X1 u2_u8_u4_U26 (.A1( u2_u8_u4_n145 ) , .A2( u2_u8_u4_n147 ) , .ZN( u2_u8_u4_n159 ) );
  OR3_X1 u2_u8_u4_U27 (.A3( u2_u8_u4_n114 ) , .A2( u2_u8_u4_n115 ) , .A1( u2_u8_u4_n116 ) , .ZN( u2_u8_u4_n136 ) );
  AOI21_X1 u2_u8_u4_U28 (.A( u2_u8_u4_n113 ) , .ZN( u2_u8_u4_n116 ) , .B2( u2_u8_u4_n173 ) , .B1( u2_u8_u4_n174 ) );
  AOI21_X1 u2_u8_u4_U29 (.ZN( u2_u8_u4_n115 ) , .B2( u2_u8_u4_n145 ) , .B1( u2_u8_u4_n146 ) , .A( u2_u8_u4_n156 ) );
  NOR2_X1 u2_u8_u4_U3 (.ZN( u2_u8_u4_n121 ) , .A1( u2_u8_u4_n181 ) , .A2( u2_u8_u4_n182 ) );
  OAI22_X1 u2_u8_u4_U30 (.ZN( u2_u8_u4_n114 ) , .A2( u2_u8_u4_n121 ) , .B1( u2_u8_u4_n160 ) , .B2( u2_u8_u4_n170 ) , .A1( u2_u8_u4_n171 ) );
  INV_X1 u2_u8_u4_U31 (.A( u2_u8_u4_n158 ) , .ZN( u2_u8_u4_n182 ) );
  INV_X1 u2_u8_u4_U32 (.ZN( u2_u8_u4_n181 ) , .A( u2_u8_u4_n96 ) );
  INV_X1 u2_u8_u4_U33 (.A( u2_u8_u4_n144 ) , .ZN( u2_u8_u4_n179 ) );
  INV_X1 u2_u8_u4_U34 (.A( u2_u8_u4_n157 ) , .ZN( u2_u8_u4_n178 ) );
  NAND2_X1 u2_u8_u4_U35 (.A2( u2_u8_u4_n154 ) , .A1( u2_u8_u4_n96 ) , .ZN( u2_u8_u4_n97 ) );
  INV_X1 u2_u8_u4_U36 (.ZN( u2_u8_u4_n186 ) , .A( u2_u8_u4_n95 ) );
  OAI221_X1 u2_u8_u4_U37 (.C1( u2_u8_u4_n134 ) , .B1( u2_u8_u4_n158 ) , .B2( u2_u8_u4_n171 ) , .C2( u2_u8_u4_n173 ) , .A( u2_u8_u4_n94 ) , .ZN( u2_u8_u4_n95 ) );
  AOI222_X1 u2_u8_u4_U38 (.B2( u2_u8_u4_n132 ) , .A1( u2_u8_u4_n138 ) , .C2( u2_u8_u4_n175 ) , .A2( u2_u8_u4_n179 ) , .C1( u2_u8_u4_n181 ) , .B1( u2_u8_u4_n185 ) , .ZN( u2_u8_u4_n94 ) );
  INV_X1 u2_u8_u4_U39 (.A( u2_u8_u4_n113 ) , .ZN( u2_u8_u4_n185 ) );
  INV_X1 u2_u8_u4_U4 (.A( u2_u8_u4_n117 ) , .ZN( u2_u8_u4_n184 ) );
  INV_X1 u2_u8_u4_U40 (.A( u2_u8_u4_n143 ) , .ZN( u2_u8_u4_n183 ) );
  NOR2_X1 u2_u8_u4_U41 (.ZN( u2_u8_u4_n138 ) , .A1( u2_u8_u4_n168 ) , .A2( u2_u8_u4_n169 ) );
  NOR2_X1 u2_u8_u4_U42 (.A1( u2_u8_u4_n150 ) , .A2( u2_u8_u4_n152 ) , .ZN( u2_u8_u4_n153 ) );
  NOR2_X1 u2_u8_u4_U43 (.A2( u2_u8_u4_n128 ) , .A1( u2_u8_u4_n138 ) , .ZN( u2_u8_u4_n156 ) );
  AOI22_X1 u2_u8_u4_U44 (.B2( u2_u8_u4_n122 ) , .A1( u2_u8_u4_n123 ) , .ZN( u2_u8_u4_n124 ) , .B1( u2_u8_u4_n128 ) , .A2( u2_u8_u4_n172 ) );
  INV_X1 u2_u8_u4_U45 (.A( u2_u8_u4_n153 ) , .ZN( u2_u8_u4_n172 ) );
  NAND2_X1 u2_u8_u4_U46 (.A2( u2_u8_u4_n120 ) , .ZN( u2_u8_u4_n123 ) , .A1( u2_u8_u4_n161 ) );
  AOI22_X1 u2_u8_u4_U47 (.B2( u2_u8_u4_n132 ) , .A2( u2_u8_u4_n133 ) , .ZN( u2_u8_u4_n140 ) , .A1( u2_u8_u4_n150 ) , .B1( u2_u8_u4_n179 ) );
  NAND2_X1 u2_u8_u4_U48 (.ZN( u2_u8_u4_n133 ) , .A2( u2_u8_u4_n146 ) , .A1( u2_u8_u4_n154 ) );
  NAND2_X1 u2_u8_u4_U49 (.A1( u2_u8_u4_n103 ) , .ZN( u2_u8_u4_n154 ) , .A2( u2_u8_u4_n98 ) );
  NOR4_X1 u2_u8_u4_U5 (.A4( u2_u8_u4_n106 ) , .A3( u2_u8_u4_n107 ) , .A2( u2_u8_u4_n108 ) , .A1( u2_u8_u4_n109 ) , .ZN( u2_u8_u4_n110 ) );
  NAND2_X1 u2_u8_u4_U50 (.A1( u2_u8_u4_n101 ) , .ZN( u2_u8_u4_n158 ) , .A2( u2_u8_u4_n99 ) );
  AOI21_X1 u2_u8_u4_U51 (.ZN( u2_u8_u4_n127 ) , .A( u2_u8_u4_n136 ) , .B2( u2_u8_u4_n150 ) , .B1( u2_u8_u4_n180 ) );
  INV_X1 u2_u8_u4_U52 (.A( u2_u8_u4_n160 ) , .ZN( u2_u8_u4_n180 ) );
  NAND2_X1 u2_u8_u4_U53 (.A2( u2_u8_u4_n104 ) , .A1( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n146 ) );
  NAND2_X1 u2_u8_u4_U54 (.A2( u2_u8_u4_n101 ) , .A1( u2_u8_u4_n102 ) , .ZN( u2_u8_u4_n160 ) );
  NAND2_X1 u2_u8_u4_U55 (.ZN( u2_u8_u4_n134 ) , .A1( u2_u8_u4_n98 ) , .A2( u2_u8_u4_n99 ) );
  NAND2_X1 u2_u8_u4_U56 (.A1( u2_u8_u4_n103 ) , .A2( u2_u8_u4_n104 ) , .ZN( u2_u8_u4_n143 ) );
  NAND2_X1 u2_u8_u4_U57 (.A2( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n145 ) , .A1( u2_u8_u4_n98 ) );
  NAND2_X1 u2_u8_u4_U58 (.A1( u2_u8_u4_n100 ) , .A2( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n120 ) );
  NAND2_X1 u2_u8_u4_U59 (.A1( u2_u8_u4_n102 ) , .A2( u2_u8_u4_n104 ) , .ZN( u2_u8_u4_n148 ) );
  AOI21_X1 u2_u8_u4_U6 (.ZN( u2_u8_u4_n106 ) , .B2( u2_u8_u4_n146 ) , .B1( u2_u8_u4_n158 ) , .A( u2_u8_u4_n170 ) );
  NAND2_X1 u2_u8_u4_U60 (.A2( u2_u8_u4_n100 ) , .A1( u2_u8_u4_n103 ) , .ZN( u2_u8_u4_n157 ) );
  INV_X1 u2_u8_u4_U61 (.A( u2_u8_u4_n150 ) , .ZN( u2_u8_u4_n173 ) );
  INV_X1 u2_u8_u4_U62 (.A( u2_u8_u4_n152 ) , .ZN( u2_u8_u4_n171 ) );
  NAND2_X1 u2_u8_u4_U63 (.A1( u2_u8_u4_n100 ) , .ZN( u2_u8_u4_n118 ) , .A2( u2_u8_u4_n99 ) );
  NAND2_X1 u2_u8_u4_U64 (.A2( u2_u8_u4_n100 ) , .A1( u2_u8_u4_n102 ) , .ZN( u2_u8_u4_n144 ) );
  NAND2_X1 u2_u8_u4_U65 (.A2( u2_u8_u4_n101 ) , .A1( u2_u8_u4_n105 ) , .ZN( u2_u8_u4_n96 ) );
  INV_X1 u2_u8_u4_U66 (.A( u2_u8_u4_n128 ) , .ZN( u2_u8_u4_n174 ) );
  NAND2_X1 u2_u8_u4_U67 (.A2( u2_u8_u4_n102 ) , .ZN( u2_u8_u4_n119 ) , .A1( u2_u8_u4_n98 ) );
  NAND2_X1 u2_u8_u4_U68 (.A2( u2_u8_u4_n101 ) , .A1( u2_u8_u4_n103 ) , .ZN( u2_u8_u4_n147 ) );
  NAND2_X1 u2_u8_u4_U69 (.A2( u2_u8_u4_n104 ) , .ZN( u2_u8_u4_n113 ) , .A1( u2_u8_u4_n99 ) );
  AOI21_X1 u2_u8_u4_U7 (.ZN( u2_u8_u4_n108 ) , .B2( u2_u8_u4_n134 ) , .B1( u2_u8_u4_n155 ) , .A( u2_u8_u4_n156 ) );
  NOR2_X1 u2_u8_u4_U70 (.A2( u2_u8_X_28 ) , .ZN( u2_u8_u4_n150 ) , .A1( u2_u8_u4_n168 ) );
  NOR2_X1 u2_u8_u4_U71 (.A2( u2_u8_X_29 ) , .ZN( u2_u8_u4_n152 ) , .A1( u2_u8_u4_n169 ) );
  NOR2_X1 u2_u8_u4_U72 (.A2( u2_u8_X_30 ) , .ZN( u2_u8_u4_n105 ) , .A1( u2_u8_u4_n176 ) );
  NOR2_X1 u2_u8_u4_U73 (.A2( u2_u8_X_26 ) , .ZN( u2_u8_u4_n100 ) , .A1( u2_u8_u4_n177 ) );
  NOR2_X1 u2_u8_u4_U74 (.A2( u2_u8_X_28 ) , .A1( u2_u8_X_29 ) , .ZN( u2_u8_u4_n128 ) );
  NOR2_X1 u2_u8_u4_U75 (.A2( u2_u8_X_27 ) , .A1( u2_u8_X_30 ) , .ZN( u2_u8_u4_n102 ) );
  NOR2_X1 u2_u8_u4_U76 (.A2( u2_u8_X_25 ) , .A1( u2_u8_X_26 ) , .ZN( u2_u8_u4_n98 ) );
  AND2_X1 u2_u8_u4_U77 (.A2( u2_u8_X_25 ) , .A1( u2_u8_X_26 ) , .ZN( u2_u8_u4_n104 ) );
  AND2_X1 u2_u8_u4_U78 (.A1( u2_u8_X_30 ) , .A2( u2_u8_u4_n176 ) , .ZN( u2_u8_u4_n99 ) );
  AND2_X1 u2_u8_u4_U79 (.A1( u2_u8_X_26 ) , .ZN( u2_u8_u4_n101 ) , .A2( u2_u8_u4_n177 ) );
  AOI21_X1 u2_u8_u4_U8 (.ZN( u2_u8_u4_n109 ) , .A( u2_u8_u4_n153 ) , .B1( u2_u8_u4_n159 ) , .B2( u2_u8_u4_n184 ) );
  AND2_X1 u2_u8_u4_U80 (.A1( u2_u8_X_27 ) , .A2( u2_u8_X_30 ) , .ZN( u2_u8_u4_n103 ) );
  INV_X1 u2_u8_u4_U81 (.A( u2_u8_X_28 ) , .ZN( u2_u8_u4_n169 ) );
  INV_X1 u2_u8_u4_U82 (.A( u2_u8_X_29 ) , .ZN( u2_u8_u4_n168 ) );
  INV_X1 u2_u8_u4_U83 (.A( u2_u8_X_25 ) , .ZN( u2_u8_u4_n177 ) );
  INV_X1 u2_u8_u4_U84 (.A( u2_u8_X_27 ) , .ZN( u2_u8_u4_n176 ) );
  NAND4_X1 u2_u8_u4_U85 (.ZN( u2_out8_25 ) , .A4( u2_u8_u4_n139 ) , .A3( u2_u8_u4_n140 ) , .A2( u2_u8_u4_n141 ) , .A1( u2_u8_u4_n142 ) );
  OAI21_X1 u2_u8_u4_U86 (.B2( u2_u8_u4_n131 ) , .ZN( u2_u8_u4_n141 ) , .A( u2_u8_u4_n175 ) , .B1( u2_u8_u4_n183 ) );
  OAI21_X1 u2_u8_u4_U87 (.A( u2_u8_u4_n128 ) , .B2( u2_u8_u4_n129 ) , .B1( u2_u8_u4_n130 ) , .ZN( u2_u8_u4_n142 ) );
  NAND4_X1 u2_u8_u4_U88 (.ZN( u2_out8_14 ) , .A4( u2_u8_u4_n124 ) , .A3( u2_u8_u4_n125 ) , .A2( u2_u8_u4_n126 ) , .A1( u2_u8_u4_n127 ) );
  AOI22_X1 u2_u8_u4_U89 (.B2( u2_u8_u4_n117 ) , .ZN( u2_u8_u4_n126 ) , .A1( u2_u8_u4_n129 ) , .B1( u2_u8_u4_n152 ) , .A2( u2_u8_u4_n175 ) );
  AOI211_X1 u2_u8_u4_U9 (.B( u2_u8_u4_n136 ) , .A( u2_u8_u4_n137 ) , .C2( u2_u8_u4_n138 ) , .ZN( u2_u8_u4_n139 ) , .C1( u2_u8_u4_n182 ) );
  AOI22_X1 u2_u8_u4_U90 (.ZN( u2_u8_u4_n125 ) , .B2( u2_u8_u4_n131 ) , .A2( u2_u8_u4_n132 ) , .B1( u2_u8_u4_n138 ) , .A1( u2_u8_u4_n178 ) );
  NAND4_X1 u2_u8_u4_U91 (.ZN( u2_out8_8 ) , .A4( u2_u8_u4_n110 ) , .A3( u2_u8_u4_n111 ) , .A2( u2_u8_u4_n112 ) , .A1( u2_u8_u4_n186 ) );
  NAND2_X1 u2_u8_u4_U92 (.ZN( u2_u8_u4_n112 ) , .A2( u2_u8_u4_n130 ) , .A1( u2_u8_u4_n150 ) );
  AOI22_X1 u2_u8_u4_U93 (.ZN( u2_u8_u4_n111 ) , .B2( u2_u8_u4_n132 ) , .A1( u2_u8_u4_n152 ) , .B1( u2_u8_u4_n178 ) , .A2( u2_u8_u4_n97 ) );
  AOI22_X1 u2_u8_u4_U94 (.B2( u2_u8_u4_n149 ) , .B1( u2_u8_u4_n150 ) , .A2( u2_u8_u4_n151 ) , .A1( u2_u8_u4_n152 ) , .ZN( u2_u8_u4_n167 ) );
  NOR4_X1 u2_u8_u4_U95 (.A4( u2_u8_u4_n162 ) , .A3( u2_u8_u4_n163 ) , .A2( u2_u8_u4_n164 ) , .A1( u2_u8_u4_n165 ) , .ZN( u2_u8_u4_n166 ) );
  NAND3_X1 u2_u8_u4_U96 (.ZN( u2_out8_3 ) , .A3( u2_u8_u4_n166 ) , .A1( u2_u8_u4_n167 ) , .A2( u2_u8_u4_n186 ) );
  NAND3_X1 u2_u8_u4_U97 (.A3( u2_u8_u4_n146 ) , .A2( u2_u8_u4_n147 ) , .A1( u2_u8_u4_n148 ) , .ZN( u2_u8_u4_n149 ) );
  NAND3_X1 u2_u8_u4_U98 (.A3( u2_u8_u4_n143 ) , .A2( u2_u8_u4_n144 ) , .A1( u2_u8_u4_n145 ) , .ZN( u2_u8_u4_n151 ) );
  NAND3_X1 u2_u8_u4_U99 (.A3( u2_u8_u4_n121 ) , .ZN( u2_u8_u4_n122 ) , .A2( u2_u8_u4_n144 ) , .A1( u2_u8_u4_n154 ) );
  XOR2_X1 u2_u9_U13 (.B( u2_K10_42 ) , .A( u2_R8_29 ) , .Z( u2_u9_X_42 ) );
  XOR2_X1 u2_u9_U14 (.B( u2_K10_41 ) , .A( u2_R8_28 ) , .Z( u2_u9_X_41 ) );
  XOR2_X1 u2_u9_U15 (.B( u2_K10_40 ) , .A( u2_R8_27 ) , .Z( u2_u9_X_40 ) );
  XOR2_X1 u2_u9_U17 (.B( u2_K10_39 ) , .A( u2_R8_26 ) , .Z( u2_u9_X_39 ) );
  XOR2_X1 u2_u9_U18 (.B( u2_K10_38 ) , .A( u2_R8_25 ) , .Z( u2_u9_X_38 ) );
  XOR2_X1 u2_u9_U19 (.B( u2_K10_37 ) , .A( u2_R8_24 ) , .Z( u2_u9_X_37 ) );
  XOR2_X1 u2_u9_U20 (.B( u2_K10_36 ) , .A( u2_R8_25 ) , .Z( u2_u9_X_36 ) );
  XOR2_X1 u2_u9_U21 (.B( u2_K10_35 ) , .A( u2_R8_24 ) , .Z( u2_u9_X_35 ) );
  XOR2_X1 u2_u9_U22 (.B( u2_K10_34 ) , .A( u2_R8_23 ) , .Z( u2_u9_X_34 ) );
  XOR2_X1 u2_u9_U23 (.B( u2_K10_33 ) , .A( u2_R8_22 ) , .Z( u2_u9_X_33 ) );
  XOR2_X1 u2_u9_U24 (.B( u2_K10_32 ) , .A( u2_R8_21 ) , .Z( u2_u9_X_32 ) );
  XOR2_X1 u2_u9_U25 (.B( u2_K10_31 ) , .A( u2_R8_20 ) , .Z( u2_u9_X_31 ) );
  NOR2_X1 u2_u9_u5_U10 (.ZN( u2_u9_u5_n135 ) , .A1( u2_u9_u5_n173 ) , .A2( u2_u9_u5_n176 ) );
  NOR3_X1 u2_u9_u5_U100 (.A3( u2_u9_u5_n141 ) , .A1( u2_u9_u5_n142 ) , .ZN( u2_u9_u5_n143 ) , .A2( u2_u9_u5_n191 ) );
  NAND4_X1 u2_u9_u5_U101 (.ZN( u2_out9_4 ) , .A4( u2_u9_u5_n112 ) , .A2( u2_u9_u5_n113 ) , .A1( u2_u9_u5_n114 ) , .A3( u2_u9_u5_n195 ) );
  AOI211_X1 u2_u9_u5_U102 (.A( u2_u9_u5_n110 ) , .C1( u2_u9_u5_n111 ) , .ZN( u2_u9_u5_n112 ) , .B( u2_u9_u5_n118 ) , .C2( u2_u9_u5_n177 ) );
  INV_X1 u2_u9_u5_U103 (.A( u2_u9_u5_n102 ) , .ZN( u2_u9_u5_n195 ) );
  NAND3_X1 u2_u9_u5_U104 (.A2( u2_u9_u5_n154 ) , .A3( u2_u9_u5_n158 ) , .A1( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n99 ) );
  INV_X1 u2_u9_u5_U11 (.A( u2_u9_u5_n121 ) , .ZN( u2_u9_u5_n177 ) );
  NOR2_X1 u2_u9_u5_U12 (.ZN( u2_u9_u5_n160 ) , .A2( u2_u9_u5_n173 ) , .A1( u2_u9_u5_n177 ) );
  INV_X1 u2_u9_u5_U13 (.A( u2_u9_u5_n150 ) , .ZN( u2_u9_u5_n174 ) );
  AOI21_X1 u2_u9_u5_U14 (.A( u2_u9_u5_n160 ) , .B2( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n162 ) , .B1( u2_u9_u5_n192 ) );
  INV_X1 u2_u9_u5_U15 (.A( u2_u9_u5_n159 ) , .ZN( u2_u9_u5_n192 ) );
  AOI21_X1 u2_u9_u5_U16 (.A( u2_u9_u5_n156 ) , .B2( u2_u9_u5_n157 ) , .B1( u2_u9_u5_n158 ) , .ZN( u2_u9_u5_n163 ) );
  AOI21_X1 u2_u9_u5_U17 (.B2( u2_u9_u5_n139 ) , .B1( u2_u9_u5_n140 ) , .ZN( u2_u9_u5_n141 ) , .A( u2_u9_u5_n150 ) );
  OAI21_X1 u2_u9_u5_U18 (.A( u2_u9_u5_n133 ) , .B2( u2_u9_u5_n134 ) , .B1( u2_u9_u5_n135 ) , .ZN( u2_u9_u5_n142 ) );
  OAI21_X1 u2_u9_u5_U19 (.ZN( u2_u9_u5_n133 ) , .B2( u2_u9_u5_n147 ) , .A( u2_u9_u5_n173 ) , .B1( u2_u9_u5_n188 ) );
  NAND2_X1 u2_u9_u5_U20 (.A2( u2_u9_u5_n119 ) , .A1( u2_u9_u5_n123 ) , .ZN( u2_u9_u5_n137 ) );
  INV_X1 u2_u9_u5_U21 (.A( u2_u9_u5_n155 ) , .ZN( u2_u9_u5_n194 ) );
  NAND2_X1 u2_u9_u5_U22 (.A1( u2_u9_u5_n121 ) , .ZN( u2_u9_u5_n132 ) , .A2( u2_u9_u5_n172 ) );
  NAND2_X1 u2_u9_u5_U23 (.A2( u2_u9_u5_n122 ) , .ZN( u2_u9_u5_n136 ) , .A1( u2_u9_u5_n154 ) );
  NAND2_X1 u2_u9_u5_U24 (.A2( u2_u9_u5_n119 ) , .A1( u2_u9_u5_n120 ) , .ZN( u2_u9_u5_n159 ) );
  INV_X1 u2_u9_u5_U25 (.A( u2_u9_u5_n156 ) , .ZN( u2_u9_u5_n175 ) );
  INV_X1 u2_u9_u5_U26 (.A( u2_u9_u5_n158 ) , .ZN( u2_u9_u5_n188 ) );
  INV_X1 u2_u9_u5_U27 (.A( u2_u9_u5_n152 ) , .ZN( u2_u9_u5_n179 ) );
  INV_X1 u2_u9_u5_U28 (.A( u2_u9_u5_n140 ) , .ZN( u2_u9_u5_n182 ) );
  INV_X1 u2_u9_u5_U29 (.A( u2_u9_u5_n151 ) , .ZN( u2_u9_u5_n183 ) );
  NOR2_X1 u2_u9_u5_U3 (.ZN( u2_u9_u5_n134 ) , .A1( u2_u9_u5_n183 ) , .A2( u2_u9_u5_n190 ) );
  INV_X1 u2_u9_u5_U30 (.A( u2_u9_u5_n123 ) , .ZN( u2_u9_u5_n185 ) );
  INV_X1 u2_u9_u5_U31 (.A( u2_u9_u5_n161 ) , .ZN( u2_u9_u5_n184 ) );
  INV_X1 u2_u9_u5_U32 (.A( u2_u9_u5_n139 ) , .ZN( u2_u9_u5_n189 ) );
  INV_X1 u2_u9_u5_U33 (.A( u2_u9_u5_n157 ) , .ZN( u2_u9_u5_n190 ) );
  INV_X1 u2_u9_u5_U34 (.A( u2_u9_u5_n120 ) , .ZN( u2_u9_u5_n193 ) );
  NAND2_X1 u2_u9_u5_U35 (.ZN( u2_u9_u5_n111 ) , .A1( u2_u9_u5_n140 ) , .A2( u2_u9_u5_n155 ) );
  NOR2_X1 u2_u9_u5_U36 (.ZN( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n170 ) , .A2( u2_u9_u5_n180 ) );
  INV_X1 u2_u9_u5_U37 (.A( u2_u9_u5_n117 ) , .ZN( u2_u9_u5_n196 ) );
  OAI221_X1 u2_u9_u5_U38 (.A( u2_u9_u5_n116 ) , .ZN( u2_u9_u5_n117 ) , .B2( u2_u9_u5_n119 ) , .C1( u2_u9_u5_n153 ) , .C2( u2_u9_u5_n158 ) , .B1( u2_u9_u5_n172 ) );
  AOI222_X1 u2_u9_u5_U39 (.ZN( u2_u9_u5_n116 ) , .B2( u2_u9_u5_n145 ) , .C1( u2_u9_u5_n148 ) , .A2( u2_u9_u5_n174 ) , .C2( u2_u9_u5_n177 ) , .B1( u2_u9_u5_n187 ) , .A1( u2_u9_u5_n193 ) );
  INV_X1 u2_u9_u5_U4 (.A( u2_u9_u5_n138 ) , .ZN( u2_u9_u5_n191 ) );
  INV_X1 u2_u9_u5_U40 (.A( u2_u9_u5_n115 ) , .ZN( u2_u9_u5_n187 ) );
  OAI221_X1 u2_u9_u5_U41 (.A( u2_u9_u5_n101 ) , .ZN( u2_u9_u5_n102 ) , .C2( u2_u9_u5_n115 ) , .C1( u2_u9_u5_n126 ) , .B1( u2_u9_u5_n134 ) , .B2( u2_u9_u5_n160 ) );
  OAI21_X1 u2_u9_u5_U42 (.ZN( u2_u9_u5_n101 ) , .B1( u2_u9_u5_n137 ) , .A( u2_u9_u5_n146 ) , .B2( u2_u9_u5_n147 ) );
  AOI22_X1 u2_u9_u5_U43 (.B2( u2_u9_u5_n131 ) , .A2( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n169 ) , .B1( u2_u9_u5_n174 ) , .A1( u2_u9_u5_n185 ) );
  NOR2_X1 u2_u9_u5_U44 (.A1( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n150 ) , .A2( u2_u9_u5_n173 ) );
  AOI21_X1 u2_u9_u5_U45 (.A( u2_u9_u5_n118 ) , .B2( u2_u9_u5_n145 ) , .ZN( u2_u9_u5_n168 ) , .B1( u2_u9_u5_n186 ) );
  INV_X1 u2_u9_u5_U46 (.A( u2_u9_u5_n122 ) , .ZN( u2_u9_u5_n186 ) );
  NOR2_X1 u2_u9_u5_U47 (.A1( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n152 ) , .A2( u2_u9_u5_n176 ) );
  NOR2_X1 u2_u9_u5_U48 (.A1( u2_u9_u5_n115 ) , .ZN( u2_u9_u5_n118 ) , .A2( u2_u9_u5_n153 ) );
  NOR2_X1 u2_u9_u5_U49 (.A2( u2_u9_u5_n145 ) , .ZN( u2_u9_u5_n156 ) , .A1( u2_u9_u5_n174 ) );
  OAI21_X1 u2_u9_u5_U5 (.B2( u2_u9_u5_n136 ) , .B1( u2_u9_u5_n137 ) , .ZN( u2_u9_u5_n138 ) , .A( u2_u9_u5_n177 ) );
  NOR2_X1 u2_u9_u5_U50 (.ZN( u2_u9_u5_n121 ) , .A2( u2_u9_u5_n145 ) , .A1( u2_u9_u5_n176 ) );
  AOI22_X1 u2_u9_u5_U51 (.ZN( u2_u9_u5_n114 ) , .A2( u2_u9_u5_n137 ) , .A1( u2_u9_u5_n145 ) , .B2( u2_u9_u5_n175 ) , .B1( u2_u9_u5_n193 ) );
  OAI211_X1 u2_u9_u5_U52 (.B( u2_u9_u5_n124 ) , .A( u2_u9_u5_n125 ) , .C2( u2_u9_u5_n126 ) , .C1( u2_u9_u5_n127 ) , .ZN( u2_u9_u5_n128 ) );
  NOR3_X1 u2_u9_u5_U53 (.ZN( u2_u9_u5_n127 ) , .A1( u2_u9_u5_n136 ) , .A3( u2_u9_u5_n148 ) , .A2( u2_u9_u5_n182 ) );
  OAI21_X1 u2_u9_u5_U54 (.ZN( u2_u9_u5_n124 ) , .A( u2_u9_u5_n177 ) , .B2( u2_u9_u5_n183 ) , .B1( u2_u9_u5_n189 ) );
  OAI21_X1 u2_u9_u5_U55 (.ZN( u2_u9_u5_n125 ) , .A( u2_u9_u5_n174 ) , .B2( u2_u9_u5_n185 ) , .B1( u2_u9_u5_n190 ) );
  AOI21_X1 u2_u9_u5_U56 (.A( u2_u9_u5_n153 ) , .B2( u2_u9_u5_n154 ) , .B1( u2_u9_u5_n155 ) , .ZN( u2_u9_u5_n164 ) );
  AOI21_X1 u2_u9_u5_U57 (.ZN( u2_u9_u5_n110 ) , .B1( u2_u9_u5_n122 ) , .B2( u2_u9_u5_n139 ) , .A( u2_u9_u5_n153 ) );
  INV_X1 u2_u9_u5_U58 (.A( u2_u9_u5_n153 ) , .ZN( u2_u9_u5_n176 ) );
  INV_X1 u2_u9_u5_U59 (.A( u2_u9_u5_n126 ) , .ZN( u2_u9_u5_n173 ) );
  AOI222_X1 u2_u9_u5_U6 (.ZN( u2_u9_u5_n113 ) , .A1( u2_u9_u5_n131 ) , .C1( u2_u9_u5_n148 ) , .B2( u2_u9_u5_n174 ) , .C2( u2_u9_u5_n178 ) , .A2( u2_u9_u5_n179 ) , .B1( u2_u9_u5_n99 ) );
  AND2_X1 u2_u9_u5_U60 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n147 ) );
  AND2_X1 u2_u9_u5_U61 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n148 ) );
  NAND2_X1 u2_u9_u5_U62 (.A1( u2_u9_u5_n105 ) , .A2( u2_u9_u5_n106 ) , .ZN( u2_u9_u5_n158 ) );
  NAND2_X1 u2_u9_u5_U63 (.A2( u2_u9_u5_n108 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n139 ) );
  NAND2_X1 u2_u9_u5_U64 (.A1( u2_u9_u5_n106 ) , .A2( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n119 ) );
  NAND2_X1 u2_u9_u5_U65 (.A2( u2_u9_u5_n103 ) , .A1( u2_u9_u5_n105 ) , .ZN( u2_u9_u5_n140 ) );
  NAND2_X1 u2_u9_u5_U66 (.A2( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n105 ) , .ZN( u2_u9_u5_n155 ) );
  NAND2_X1 u2_u9_u5_U67 (.A2( u2_u9_u5_n106 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n122 ) );
  NAND2_X1 u2_u9_u5_U68 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n106 ) , .ZN( u2_u9_u5_n115 ) );
  NAND2_X1 u2_u9_u5_U69 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n103 ) , .ZN( u2_u9_u5_n161 ) );
  INV_X1 u2_u9_u5_U7 (.A( u2_u9_u5_n135 ) , .ZN( u2_u9_u5_n178 ) );
  NAND2_X1 u2_u9_u5_U70 (.A1( u2_u9_u5_n105 ) , .A2( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n154 ) );
  INV_X1 u2_u9_u5_U71 (.A( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n172 ) );
  NAND2_X1 u2_u9_u5_U72 (.A1( u2_u9_u5_n103 ) , .A2( u2_u9_u5_n108 ) , .ZN( u2_u9_u5_n123 ) );
  NAND2_X1 u2_u9_u5_U73 (.A2( u2_u9_u5_n103 ) , .A1( u2_u9_u5_n107 ) , .ZN( u2_u9_u5_n151 ) );
  NAND2_X1 u2_u9_u5_U74 (.A2( u2_u9_u5_n107 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n120 ) );
  NAND2_X1 u2_u9_u5_U75 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n109 ) , .ZN( u2_u9_u5_n157 ) );
  AND2_X1 u2_u9_u5_U76 (.A2( u2_u9_u5_n100 ) , .A1( u2_u9_u5_n104 ) , .ZN( u2_u9_u5_n131 ) );
  NOR2_X1 u2_u9_u5_U77 (.A2( u2_u9_X_34 ) , .A1( u2_u9_X_35 ) , .ZN( u2_u9_u5_n145 ) );
  NOR2_X1 u2_u9_u5_U78 (.A2( u2_u9_X_34 ) , .ZN( u2_u9_u5_n146 ) , .A1( u2_u9_u5_n171 ) );
  NOR2_X1 u2_u9_u5_U79 (.A2( u2_u9_X_31 ) , .A1( u2_u9_X_32 ) , .ZN( u2_u9_u5_n103 ) );
  OAI22_X1 u2_u9_u5_U8 (.B2( u2_u9_u5_n149 ) , .B1( u2_u9_u5_n150 ) , .A2( u2_u9_u5_n151 ) , .A1( u2_u9_u5_n152 ) , .ZN( u2_u9_u5_n165 ) );
  NOR2_X1 u2_u9_u5_U80 (.A2( u2_u9_X_36 ) , .ZN( u2_u9_u5_n105 ) , .A1( u2_u9_u5_n180 ) );
  NOR2_X1 u2_u9_u5_U81 (.A2( u2_u9_X_33 ) , .ZN( u2_u9_u5_n108 ) , .A1( u2_u9_u5_n170 ) );
  NOR2_X1 u2_u9_u5_U82 (.A2( u2_u9_X_33 ) , .A1( u2_u9_X_36 ) , .ZN( u2_u9_u5_n107 ) );
  NOR2_X1 u2_u9_u5_U83 (.A2( u2_u9_X_31 ) , .ZN( u2_u9_u5_n104 ) , .A1( u2_u9_u5_n181 ) );
  NAND2_X1 u2_u9_u5_U84 (.A2( u2_u9_X_34 ) , .A1( u2_u9_X_35 ) , .ZN( u2_u9_u5_n153 ) );
  NAND2_X1 u2_u9_u5_U85 (.A1( u2_u9_X_34 ) , .ZN( u2_u9_u5_n126 ) , .A2( u2_u9_u5_n171 ) );
  AND2_X1 u2_u9_u5_U86 (.A1( u2_u9_X_31 ) , .A2( u2_u9_X_32 ) , .ZN( u2_u9_u5_n106 ) );
  AND2_X1 u2_u9_u5_U87 (.A1( u2_u9_X_31 ) , .ZN( u2_u9_u5_n109 ) , .A2( u2_u9_u5_n181 ) );
  INV_X1 u2_u9_u5_U88 (.A( u2_u9_X_33 ) , .ZN( u2_u9_u5_n180 ) );
  INV_X1 u2_u9_u5_U89 (.A( u2_u9_X_35 ) , .ZN( u2_u9_u5_n171 ) );
  NOR3_X1 u2_u9_u5_U9 (.A2( u2_u9_u5_n147 ) , .A1( u2_u9_u5_n148 ) , .ZN( u2_u9_u5_n149 ) , .A3( u2_u9_u5_n194 ) );
  INV_X1 u2_u9_u5_U90 (.A( u2_u9_X_36 ) , .ZN( u2_u9_u5_n170 ) );
  INV_X1 u2_u9_u5_U91 (.A( u2_u9_X_32 ) , .ZN( u2_u9_u5_n181 ) );
  NAND4_X1 u2_u9_u5_U92 (.ZN( u2_out9_29 ) , .A4( u2_u9_u5_n129 ) , .A3( u2_u9_u5_n130 ) , .A2( u2_u9_u5_n168 ) , .A1( u2_u9_u5_n196 ) );
  AOI221_X1 u2_u9_u5_U93 (.A( u2_u9_u5_n128 ) , .ZN( u2_u9_u5_n129 ) , .C2( u2_u9_u5_n132 ) , .B2( u2_u9_u5_n159 ) , .B1( u2_u9_u5_n176 ) , .C1( u2_u9_u5_n184 ) );
  AOI222_X1 u2_u9_u5_U94 (.ZN( u2_u9_u5_n130 ) , .A2( u2_u9_u5_n146 ) , .B1( u2_u9_u5_n147 ) , .C2( u2_u9_u5_n175 ) , .B2( u2_u9_u5_n179 ) , .A1( u2_u9_u5_n188 ) , .C1( u2_u9_u5_n194 ) );
  NAND4_X1 u2_u9_u5_U95 (.ZN( u2_out9_19 ) , .A4( u2_u9_u5_n166 ) , .A3( u2_u9_u5_n167 ) , .A2( u2_u9_u5_n168 ) , .A1( u2_u9_u5_n169 ) );
  AOI22_X1 u2_u9_u5_U96 (.B2( u2_u9_u5_n145 ) , .A2( u2_u9_u5_n146 ) , .ZN( u2_u9_u5_n167 ) , .B1( u2_u9_u5_n182 ) , .A1( u2_u9_u5_n189 ) );
  NOR4_X1 u2_u9_u5_U97 (.A4( u2_u9_u5_n162 ) , .A3( u2_u9_u5_n163 ) , .A2( u2_u9_u5_n164 ) , .A1( u2_u9_u5_n165 ) , .ZN( u2_u9_u5_n166 ) );
  NAND4_X1 u2_u9_u5_U98 (.ZN( u2_out9_11 ) , .A4( u2_u9_u5_n143 ) , .A3( u2_u9_u5_n144 ) , .A2( u2_u9_u5_n169 ) , .A1( u2_u9_u5_n196 ) );
  AOI22_X1 u2_u9_u5_U99 (.A2( u2_u9_u5_n132 ) , .ZN( u2_u9_u5_n144 ) , .B2( u2_u9_u5_n145 ) , .B1( u2_u9_u5_n184 ) , .A1( u2_u9_u5_n194 ) );
  AOI22_X1 u2_u9_u6_U10 (.A2( u2_u9_u6_n151 ) , .B2( u2_u9_u6_n161 ) , .A1( u2_u9_u6_n167 ) , .B1( u2_u9_u6_n170 ) , .ZN( u2_u9_u6_n89 ) );
  AOI21_X1 u2_u9_u6_U11 (.B1( u2_u9_u6_n107 ) , .B2( u2_u9_u6_n132 ) , .A( u2_u9_u6_n158 ) , .ZN( u2_u9_u6_n88 ) );
  AOI21_X1 u2_u9_u6_U12 (.B2( u2_u9_u6_n147 ) , .B1( u2_u9_u6_n148 ) , .ZN( u2_u9_u6_n149 ) , .A( u2_u9_u6_n158 ) );
  AOI21_X1 u2_u9_u6_U13 (.ZN( u2_u9_u6_n106 ) , .A( u2_u9_u6_n142 ) , .B2( u2_u9_u6_n159 ) , .B1( u2_u9_u6_n164 ) );
  INV_X1 u2_u9_u6_U14 (.A( u2_u9_u6_n155 ) , .ZN( u2_u9_u6_n161 ) );
  INV_X1 u2_u9_u6_U15 (.A( u2_u9_u6_n128 ) , .ZN( u2_u9_u6_n164 ) );
  NAND2_X1 u2_u9_u6_U16 (.ZN( u2_u9_u6_n110 ) , .A1( u2_u9_u6_n122 ) , .A2( u2_u9_u6_n129 ) );
  NAND2_X1 u2_u9_u6_U17 (.ZN( u2_u9_u6_n124 ) , .A2( u2_u9_u6_n146 ) , .A1( u2_u9_u6_n148 ) );
  INV_X1 u2_u9_u6_U18 (.A( u2_u9_u6_n132 ) , .ZN( u2_u9_u6_n171 ) );
  AND2_X1 u2_u9_u6_U19 (.A1( u2_u9_u6_n100 ) , .ZN( u2_u9_u6_n130 ) , .A2( u2_u9_u6_n147 ) );
  INV_X1 u2_u9_u6_U20 (.A( u2_u9_u6_n127 ) , .ZN( u2_u9_u6_n173 ) );
  INV_X1 u2_u9_u6_U21 (.A( u2_u9_u6_n121 ) , .ZN( u2_u9_u6_n167 ) );
  INV_X1 u2_u9_u6_U22 (.A( u2_u9_u6_n100 ) , .ZN( u2_u9_u6_n169 ) );
  INV_X1 u2_u9_u6_U23 (.A( u2_u9_u6_n123 ) , .ZN( u2_u9_u6_n170 ) );
  INV_X1 u2_u9_u6_U24 (.A( u2_u9_u6_n113 ) , .ZN( u2_u9_u6_n168 ) );
  AND2_X1 u2_u9_u6_U25 (.A1( u2_u9_u6_n107 ) , .A2( u2_u9_u6_n119 ) , .ZN( u2_u9_u6_n133 ) );
  AND2_X1 u2_u9_u6_U26 (.A2( u2_u9_u6_n121 ) , .A1( u2_u9_u6_n122 ) , .ZN( u2_u9_u6_n131 ) );
  AND3_X1 u2_u9_u6_U27 (.ZN( u2_u9_u6_n120 ) , .A2( u2_u9_u6_n127 ) , .A1( u2_u9_u6_n132 ) , .A3( u2_u9_u6_n145 ) );
  INV_X1 u2_u9_u6_U28 (.A( u2_u9_u6_n146 ) , .ZN( u2_u9_u6_n163 ) );
  AOI222_X1 u2_u9_u6_U29 (.ZN( u2_u9_u6_n114 ) , .A1( u2_u9_u6_n118 ) , .A2( u2_u9_u6_n126 ) , .B2( u2_u9_u6_n151 ) , .C2( u2_u9_u6_n159 ) , .C1( u2_u9_u6_n168 ) , .B1( u2_u9_u6_n169 ) );
  INV_X1 u2_u9_u6_U3 (.A( u2_u9_u6_n110 ) , .ZN( u2_u9_u6_n166 ) );
  NOR2_X1 u2_u9_u6_U30 (.A1( u2_u9_u6_n162 ) , .A2( u2_u9_u6_n165 ) , .ZN( u2_u9_u6_n98 ) );
  NAND2_X1 u2_u9_u6_U31 (.A1( u2_u9_u6_n144 ) , .ZN( u2_u9_u6_n151 ) , .A2( u2_u9_u6_n158 ) );
  NAND2_X1 u2_u9_u6_U32 (.ZN( u2_u9_u6_n132 ) , .A1( u2_u9_u6_n91 ) , .A2( u2_u9_u6_n97 ) );
  AOI22_X1 u2_u9_u6_U33 (.B2( u2_u9_u6_n110 ) , .B1( u2_u9_u6_n111 ) , .A1( u2_u9_u6_n112 ) , .ZN( u2_u9_u6_n115 ) , .A2( u2_u9_u6_n161 ) );
  NAND4_X1 u2_u9_u6_U34 (.A3( u2_u9_u6_n109 ) , .ZN( u2_u9_u6_n112 ) , .A4( u2_u9_u6_n132 ) , .A2( u2_u9_u6_n147 ) , .A1( u2_u9_u6_n166 ) );
  NOR2_X1 u2_u9_u6_U35 (.ZN( u2_u9_u6_n109 ) , .A1( u2_u9_u6_n170 ) , .A2( u2_u9_u6_n173 ) );
  NOR2_X1 u2_u9_u6_U36 (.A2( u2_u9_u6_n126 ) , .ZN( u2_u9_u6_n155 ) , .A1( u2_u9_u6_n160 ) );
  NAND2_X1 u2_u9_u6_U37 (.ZN( u2_u9_u6_n146 ) , .A2( u2_u9_u6_n94 ) , .A1( u2_u9_u6_n99 ) );
  AOI21_X1 u2_u9_u6_U38 (.A( u2_u9_u6_n144 ) , .B2( u2_u9_u6_n145 ) , .B1( u2_u9_u6_n146 ) , .ZN( u2_u9_u6_n150 ) );
  AOI211_X1 u2_u9_u6_U39 (.B( u2_u9_u6_n134 ) , .A( u2_u9_u6_n135 ) , .C1( u2_u9_u6_n136 ) , .ZN( u2_u9_u6_n137 ) , .C2( u2_u9_u6_n151 ) );
  INV_X1 u2_u9_u6_U4 (.A( u2_u9_u6_n142 ) , .ZN( u2_u9_u6_n174 ) );
  NAND4_X1 u2_u9_u6_U40 (.A4( u2_u9_u6_n127 ) , .A3( u2_u9_u6_n128 ) , .A2( u2_u9_u6_n129 ) , .A1( u2_u9_u6_n130 ) , .ZN( u2_u9_u6_n136 ) );
  AOI21_X1 u2_u9_u6_U41 (.B2( u2_u9_u6_n132 ) , .B1( u2_u9_u6_n133 ) , .ZN( u2_u9_u6_n134 ) , .A( u2_u9_u6_n158 ) );
  AOI21_X1 u2_u9_u6_U42 (.B1( u2_u9_u6_n131 ) , .ZN( u2_u9_u6_n135 ) , .A( u2_u9_u6_n144 ) , .B2( u2_u9_u6_n146 ) );
  INV_X1 u2_u9_u6_U43 (.A( u2_u9_u6_n111 ) , .ZN( u2_u9_u6_n158 ) );
  NAND2_X1 u2_u9_u6_U44 (.ZN( u2_u9_u6_n127 ) , .A1( u2_u9_u6_n91 ) , .A2( u2_u9_u6_n92 ) );
  NAND2_X1 u2_u9_u6_U45 (.ZN( u2_u9_u6_n129 ) , .A2( u2_u9_u6_n95 ) , .A1( u2_u9_u6_n96 ) );
  INV_X1 u2_u9_u6_U46 (.A( u2_u9_u6_n144 ) , .ZN( u2_u9_u6_n159 ) );
  NAND2_X1 u2_u9_u6_U47 (.ZN( u2_u9_u6_n145 ) , .A2( u2_u9_u6_n97 ) , .A1( u2_u9_u6_n98 ) );
  NAND2_X1 u2_u9_u6_U48 (.ZN( u2_u9_u6_n148 ) , .A2( u2_u9_u6_n92 ) , .A1( u2_u9_u6_n94 ) );
  NAND2_X1 u2_u9_u6_U49 (.ZN( u2_u9_u6_n108 ) , .A2( u2_u9_u6_n139 ) , .A1( u2_u9_u6_n144 ) );
  NAND2_X1 u2_u9_u6_U5 (.A2( u2_u9_u6_n143 ) , .ZN( u2_u9_u6_n152 ) , .A1( u2_u9_u6_n166 ) );
  NAND2_X1 u2_u9_u6_U50 (.ZN( u2_u9_u6_n121 ) , .A2( u2_u9_u6_n95 ) , .A1( u2_u9_u6_n97 ) );
  NAND2_X1 u2_u9_u6_U51 (.ZN( u2_u9_u6_n107 ) , .A2( u2_u9_u6_n92 ) , .A1( u2_u9_u6_n95 ) );
  AND2_X1 u2_u9_u6_U52 (.ZN( u2_u9_u6_n118 ) , .A2( u2_u9_u6_n91 ) , .A1( u2_u9_u6_n99 ) );
  NAND2_X1 u2_u9_u6_U53 (.ZN( u2_u9_u6_n147 ) , .A2( u2_u9_u6_n98 ) , .A1( u2_u9_u6_n99 ) );
  NAND2_X1 u2_u9_u6_U54 (.ZN( u2_u9_u6_n128 ) , .A1( u2_u9_u6_n94 ) , .A2( u2_u9_u6_n96 ) );
  NAND2_X1 u2_u9_u6_U55 (.ZN( u2_u9_u6_n119 ) , .A2( u2_u9_u6_n95 ) , .A1( u2_u9_u6_n99 ) );
  NAND2_X1 u2_u9_u6_U56 (.ZN( u2_u9_u6_n123 ) , .A2( u2_u9_u6_n91 ) , .A1( u2_u9_u6_n96 ) );
  NAND2_X1 u2_u9_u6_U57 (.ZN( u2_u9_u6_n100 ) , .A2( u2_u9_u6_n92 ) , .A1( u2_u9_u6_n98 ) );
  NAND2_X1 u2_u9_u6_U58 (.ZN( u2_u9_u6_n122 ) , .A1( u2_u9_u6_n94 ) , .A2( u2_u9_u6_n97 ) );
  INV_X1 u2_u9_u6_U59 (.A( u2_u9_u6_n139 ) , .ZN( u2_u9_u6_n160 ) );
  AOI22_X1 u2_u9_u6_U6 (.B2( u2_u9_u6_n101 ) , .A1( u2_u9_u6_n102 ) , .ZN( u2_u9_u6_n103 ) , .B1( u2_u9_u6_n160 ) , .A2( u2_u9_u6_n161 ) );
  NAND2_X1 u2_u9_u6_U60 (.ZN( u2_u9_u6_n113 ) , .A1( u2_u9_u6_n96 ) , .A2( u2_u9_u6_n98 ) );
  NOR2_X1 u2_u9_u6_U61 (.A2( u2_u9_X_40 ) , .A1( u2_u9_X_41 ) , .ZN( u2_u9_u6_n126 ) );
  NOR2_X1 u2_u9_u6_U62 (.A2( u2_u9_X_39 ) , .A1( u2_u9_X_42 ) , .ZN( u2_u9_u6_n92 ) );
  NOR2_X1 u2_u9_u6_U63 (.A2( u2_u9_X_39 ) , .A1( u2_u9_u6_n156 ) , .ZN( u2_u9_u6_n97 ) );
  NOR2_X1 u2_u9_u6_U64 (.A2( u2_u9_X_38 ) , .A1( u2_u9_u6_n165 ) , .ZN( u2_u9_u6_n95 ) );
  NOR2_X1 u2_u9_u6_U65 (.A2( u2_u9_X_41 ) , .ZN( u2_u9_u6_n111 ) , .A1( u2_u9_u6_n157 ) );
  NOR2_X1 u2_u9_u6_U66 (.A2( u2_u9_X_37 ) , .A1( u2_u9_u6_n162 ) , .ZN( u2_u9_u6_n94 ) );
  NOR2_X1 u2_u9_u6_U67 (.A2( u2_u9_X_37 ) , .A1( u2_u9_X_38 ) , .ZN( u2_u9_u6_n91 ) );
  NAND2_X1 u2_u9_u6_U68 (.A1( u2_u9_X_41 ) , .ZN( u2_u9_u6_n144 ) , .A2( u2_u9_u6_n157 ) );
  NAND2_X1 u2_u9_u6_U69 (.A2( u2_u9_X_40 ) , .A1( u2_u9_X_41 ) , .ZN( u2_u9_u6_n139 ) );
  NOR2_X1 u2_u9_u6_U7 (.A1( u2_u9_u6_n118 ) , .ZN( u2_u9_u6_n143 ) , .A2( u2_u9_u6_n168 ) );
  AND2_X1 u2_u9_u6_U70 (.A1( u2_u9_X_39 ) , .A2( u2_u9_u6_n156 ) , .ZN( u2_u9_u6_n96 ) );
  AND2_X1 u2_u9_u6_U71 (.A1( u2_u9_X_39 ) , .A2( u2_u9_X_42 ) , .ZN( u2_u9_u6_n99 ) );
  INV_X1 u2_u9_u6_U72 (.A( u2_u9_X_40 ) , .ZN( u2_u9_u6_n157 ) );
  INV_X1 u2_u9_u6_U73 (.A( u2_u9_X_37 ) , .ZN( u2_u9_u6_n165 ) );
  INV_X1 u2_u9_u6_U74 (.A( u2_u9_X_38 ) , .ZN( u2_u9_u6_n162 ) );
  INV_X1 u2_u9_u6_U75 (.A( u2_u9_X_42 ) , .ZN( u2_u9_u6_n156 ) );
  NAND4_X1 u2_u9_u6_U76 (.ZN( u2_out9_32 ) , .A4( u2_u9_u6_n103 ) , .A3( u2_u9_u6_n104 ) , .A2( u2_u9_u6_n105 ) , .A1( u2_u9_u6_n106 ) );
  AOI22_X1 u2_u9_u6_U77 (.ZN( u2_u9_u6_n105 ) , .A2( u2_u9_u6_n108 ) , .A1( u2_u9_u6_n118 ) , .B2( u2_u9_u6_n126 ) , .B1( u2_u9_u6_n171 ) );
  AOI22_X1 u2_u9_u6_U78 (.ZN( u2_u9_u6_n104 ) , .A1( u2_u9_u6_n111 ) , .B1( u2_u9_u6_n124 ) , .B2( u2_u9_u6_n151 ) , .A2( u2_u9_u6_n93 ) );
  NAND4_X1 u2_u9_u6_U79 (.ZN( u2_out9_12 ) , .A4( u2_u9_u6_n114 ) , .A3( u2_u9_u6_n115 ) , .A2( u2_u9_u6_n116 ) , .A1( u2_u9_u6_n117 ) );
  OAI21_X1 u2_u9_u6_U8 (.A( u2_u9_u6_n159 ) , .B1( u2_u9_u6_n169 ) , .B2( u2_u9_u6_n173 ) , .ZN( u2_u9_u6_n90 ) );
  OAI22_X1 u2_u9_u6_U80 (.B2( u2_u9_u6_n111 ) , .ZN( u2_u9_u6_n116 ) , .B1( u2_u9_u6_n126 ) , .A2( u2_u9_u6_n164 ) , .A1( u2_u9_u6_n167 ) );
  OAI21_X1 u2_u9_u6_U81 (.A( u2_u9_u6_n108 ) , .ZN( u2_u9_u6_n117 ) , .B2( u2_u9_u6_n141 ) , .B1( u2_u9_u6_n163 ) );
  OAI211_X1 u2_u9_u6_U82 (.ZN( u2_out9_7 ) , .B( u2_u9_u6_n153 ) , .C2( u2_u9_u6_n154 ) , .C1( u2_u9_u6_n155 ) , .A( u2_u9_u6_n174 ) );
  NOR3_X1 u2_u9_u6_U83 (.A1( u2_u9_u6_n141 ) , .ZN( u2_u9_u6_n154 ) , .A3( u2_u9_u6_n164 ) , .A2( u2_u9_u6_n171 ) );
  AOI211_X1 u2_u9_u6_U84 (.B( u2_u9_u6_n149 ) , .A( u2_u9_u6_n150 ) , .C2( u2_u9_u6_n151 ) , .C1( u2_u9_u6_n152 ) , .ZN( u2_u9_u6_n153 ) );
  OAI211_X1 u2_u9_u6_U85 (.ZN( u2_out9_22 ) , .B( u2_u9_u6_n137 ) , .A( u2_u9_u6_n138 ) , .C2( u2_u9_u6_n139 ) , .C1( u2_u9_u6_n140 ) );
  AOI22_X1 u2_u9_u6_U86 (.B1( u2_u9_u6_n124 ) , .A2( u2_u9_u6_n125 ) , .A1( u2_u9_u6_n126 ) , .ZN( u2_u9_u6_n138 ) , .B2( u2_u9_u6_n161 ) );
  AND4_X1 u2_u9_u6_U87 (.A3( u2_u9_u6_n119 ) , .A1( u2_u9_u6_n120 ) , .A4( u2_u9_u6_n129 ) , .ZN( u2_u9_u6_n140 ) , .A2( u2_u9_u6_n143 ) );
  NAND3_X1 u2_u9_u6_U88 (.A2( u2_u9_u6_n123 ) , .ZN( u2_u9_u6_n125 ) , .A1( u2_u9_u6_n130 ) , .A3( u2_u9_u6_n131 ) );
  NAND3_X1 u2_u9_u6_U89 (.A3( u2_u9_u6_n133 ) , .ZN( u2_u9_u6_n141 ) , .A1( u2_u9_u6_n145 ) , .A2( u2_u9_u6_n148 ) );
  INV_X1 u2_u9_u6_U9 (.ZN( u2_u9_u6_n172 ) , .A( u2_u9_u6_n88 ) );
  NAND3_X1 u2_u9_u6_U90 (.ZN( u2_u9_u6_n101 ) , .A3( u2_u9_u6_n107 ) , .A2( u2_u9_u6_n121 ) , .A1( u2_u9_u6_n127 ) );
  NAND3_X1 u2_u9_u6_U91 (.ZN( u2_u9_u6_n102 ) , .A3( u2_u9_u6_n130 ) , .A2( u2_u9_u6_n145 ) , .A1( u2_u9_u6_n166 ) );
  NAND3_X1 u2_u9_u6_U92 (.A3( u2_u9_u6_n113 ) , .A1( u2_u9_u6_n119 ) , .A2( u2_u9_u6_n123 ) , .ZN( u2_u9_u6_n93 ) );
  NAND3_X1 u2_u9_u6_U93 (.ZN( u2_u9_u6_n142 ) , .A2( u2_u9_u6_n172 ) , .A3( u2_u9_u6_n89 ) , .A1( u2_u9_u6_n90 ) );
  OAI21_X1 u2_uk_U1003 (.ZN( u2_K12_7 ) , .B1( u2_uk_n11 ) , .B2( u2_uk_n1720 ) , .A( u2_uk_n520 ) );
  OAI21_X1 u2_uk_U1011 (.ZN( u2_K14_44 ) , .B2( u2_uk_n1777 ) , .B1( u2_uk_n238 ) , .A( u2_uk_n717 ) );
  NAND2_X1 u2_uk_U1012 (.A1( u2_uk_K_r12_15 ) , .A2( u2_uk_n214 ) , .ZN( u2_uk_n717 ) );
  INV_X1 u2_uk_U1043 (.A( u2_key_r_9 ) , .ZN( u2_uk_n1149 ) );
  INV_X1 u2_uk_U1044 (.A( u2_key_r_7 ) , .ZN( u2_uk_n1147 ) );
  INV_X1 u2_uk_U1047 (.A( u2_key_r_23 ) , .ZN( u2_uk_n1158 ) );
  INV_X1 u2_uk_U1049 (.A( u2_key_r_30 ) , .ZN( u2_uk_n1165 ) );
  INV_X1 u2_uk_U1050 (.A( u2_key_r_47 ) , .ZN( u2_uk_n1179 ) );
  INV_X1 u2_uk_U1055 (.A( u2_key_r_37 ) , .ZN( u2_uk_n1171 ) );
  INV_X1 u2_uk_U1056 (.A( u2_key_r_52 ) , .ZN( u2_uk_n1183 ) );
  INV_X1 u2_uk_U1057 (.A( u2_key_r_0 ) , .ZN( u2_uk_n1142 ) );
  INV_X1 u2_uk_U1058 (.A( u2_key_r_16 ) , .ZN( u2_uk_n1152 ) );
  OAI22_X1 u2_uk_U106 (.ZN( u2_K10_41 ) , .A2( u2_uk_n1594 ) , .B2( u2_uk_n1622 ) , .B1( u2_uk_n17 ) , .A1( u2_uk_n231 ) );
  INV_X1 u2_uk_U1061 (.A( u2_key_r_2 ) , .ZN( u2_uk_n1144 ) );
  OAI21_X1 u2_uk_U1068 (.ZN( u2_K8_14 ) , .A( u2_uk_n1099 ) , .B2( u2_uk_n1529 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U1069 (.A1( u2_uk_K_r6_34 ) , .ZN( u2_uk_n1099 ) , .A2( u2_uk_n155 ) );
  INV_X1 u2_uk_U1080 (.A( u2_key_r_40 ) , .ZN( u2_uk_n1174 ) );
  INV_X1 u2_uk_U1088 (.ZN( u2_K8_3 ) , .A( u2_uk_n1110 ) );
  AOI22_X1 u2_uk_U1089 (.B2( u2_uk_K_r6_10 ) , .A2( u2_uk_K_r6_3 ) , .ZN( u2_uk_n1110 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n162 ) );
  INV_X1 u2_uk_U1092 (.ZN( u2_K1_41 ) , .A( u2_uk_n985 ) );
  AOI22_X1 u2_uk_U1093 (.B2( u2_key_r_35 ) , .A2( u2_key_r_42 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n60 ) , .ZN( u2_uk_n985 ) );
  INV_X1 u2_uk_U1100 (.ZN( u2_K1_20 ) , .A( u2_uk_n973 ) );
  AOI22_X1 u2_uk_U1101 (.B2( u2_key_r_48 ) , .A2( u2_key_r_55 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n63 ) , .ZN( u2_uk_n973 ) );
  INV_X1 u2_uk_U1102 (.ZN( u2_K2_32 ) , .A( u2_uk_n999 ) );
  AOI22_X1 u2_uk_U1103 (.B2( u2_uk_K_r0_15 ) , .A2( u2_uk_K_r0_36 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n155 ) , .ZN( u2_uk_n999 ) );
  INV_X1 u2_uk_U1112 (.ZN( u2_K9_20 ) , .A( u2_uk_n1126 ) );
  AOI22_X1 u2_uk_U1113 (.B2( u2_uk_K_r7_32 ) , .A2( u2_uk_K_r7_39 ) , .ZN( u2_uk_n1126 ) , .A1( u2_uk_n162 ) , .B1( u2_uk_n63 ) );
  INV_X1 u2_uk_U1114 (.ZN( u2_K5_20 ) , .A( u2_uk_n1043 ) );
  INV_X1 u2_uk_U1118 (.ZN( u2_K1_32 ) , .A( u2_uk_n980 ) );
  AOI22_X1 u2_uk_U1119 (.B2( u2_key_r_22 ) , .A2( u2_key_r_29 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n980 ) );
  INV_X1 u2_uk_U1136 (.ZN( u2_K8_15 ) , .A( u2_uk_n1100 ) );
  INV_X1 u2_uk_U1145 (.ZN( u2_K12_1 ) , .A( u2_uk_n421 ) );
  OAI22_X1 u2_uk_U1150 (.ZN( u2_K1_23 ) , .B2( u2_uk_n1167 ) , .A2( u2_uk_n1174 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n238 ) );
  INV_X1 u2_uk_U1151 (.A( u2_key_r_33 ) , .ZN( u2_uk_n1167 ) );
  OAI21_X1 u2_uk_U126 (.ZN( u2_K5_15 ) , .A( u2_uk_n1042 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1379 ) );
  INV_X1 u2_uk_U13 (.A( u2_uk_n182 ) , .ZN( u2_uk_n92 ) );
  INV_X1 u2_uk_U151 (.ZN( u2_K9_19 ) , .A( u2_uk_n1124 ) );
  AOI22_X1 u2_uk_U152 (.B1( u2_uk_K_r7_13 ) , .A2( u2_uk_K_r7_20 ) , .B2( u2_uk_n10 ) , .ZN( u2_uk_n1124 ) , .A1( u2_uk_n162 ) );
  OAI22_X1 u2_uk_U161 (.ZN( u2_K5_30 ) , .B2( u2_uk_n1378 ) , .A2( u2_uk_n1395 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n93 ) );
  OAI21_X1 u2_uk_U200 (.ZN( u2_K1_30 ) , .B1( u2_uk_n100 ) , .B2( u2_uk_n1183 ) , .A( u2_uk_n979 ) );
  OAI21_X1 u2_uk_U202 (.ZN( u2_K9_30 ) , .B1( u2_uk_n109 ) , .A( u2_uk_n1131 ) , .B2( u2_uk_n1570 ) );
  OAI22_X1 u2_uk_U211 (.ZN( u2_K1_31 ) , .A2( u2_uk_n1147 ) , .B2( u2_uk_n1151 ) , .A1( u2_uk_n208 ) , .B1( u2_uk_n31 ) );
  INV_X1 u2_uk_U212 (.A( u2_key_r_14 ) , .ZN( u2_uk_n1151 ) );
  OAI22_X1 u2_uk_U219 (.ZN( u2_K2_31 ) , .B2( u2_uk_n1230 ) , .A2( u2_uk_n1245 ) , .B1( u2_uk_n223 ) , .A1( u2_uk_n92 ) );
  INV_X1 u2_uk_U222 (.ZN( u2_K10_39 ) , .A( u2_uk_n305 ) );
  AOI22_X1 u2_uk_U223 (.B2( u2_uk_K_r8_44 ) , .A2( u2_uk_K_r8_52 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n187 ) , .ZN( u2_uk_n305 ) );
  OAI21_X1 u2_uk_U225 (.ZN( u2_K10_31 ) , .B2( u2_uk_n1615 ) , .B1( u2_uk_n164 ) , .A( u2_uk_n291 ) );
  NAND2_X1 u2_uk_U226 (.A1( u2_uk_K_r8_16 ) , .A2( u2_uk_n155 ) , .ZN( u2_uk_n291 ) );
  BUF_X1 u2_uk_U23 (.Z( u2_uk_n155 ) , .A( u2_uk_n214 ) );
  OAI21_X1 u2_uk_U232 (.ZN( u2_K1_39 ) , .B2( u2_uk_n1157 ) , .B1( u2_uk_n63 ) , .A( u2_uk_n984 ) );
  INV_X1 u2_uk_U234 (.A( u2_key_r_22 ) , .ZN( u2_uk_n1157 ) );
  INV_X1 u2_uk_U247 (.ZN( u2_K1_48 ) , .A( u2_uk_n989 ) );
  AOI22_X1 u2_uk_U248 (.B2( u2_key_r_21 ) , .A2( u2_key_r_28 ) , .B1( u2_uk_n100 ) , .A1( u2_uk_n217 ) , .ZN( u2_uk_n989 ) );
  OAI22_X1 u2_uk_U252 (.ZN( u2_K14_48 ) , .B2( u2_uk_n1768 ) , .A2( u2_uk_n1806 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n92 ) );
  BUF_X1 u2_uk_U26 (.Z( u2_uk_n148 ) , .A( u2_uk_n217 ) );
  INV_X1 u2_uk_U298 (.ZN( u2_K1_26 ) , .A( u2_uk_n976 ) );
  AOI22_X1 u2_uk_U299 (.B2( u2_key_r_31 ) , .A2( u2_key_r_51 ) , .A1( u2_uk_n118 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n976 ) );
  INV_X1 u2_uk_U301 (.ZN( u2_K9_26 ) , .A( u2_uk_n1128 ) );
  BUF_X1 u2_uk_U33 (.Z( u2_uk_n182 ) , .A( u2_uk_n208 ) );
  INV_X1 u2_uk_U338 (.ZN( u2_K12_4 ) , .A( u2_uk_n515 ) );
  AOI22_X1 u2_uk_U339 (.B2( u2_uk_K_r10_27 ) , .A2( u2_uk_K_r10_4 ) , .B1( u2_uk_n10 ) , .A1( u2_uk_n238 ) , .ZN( u2_uk_n515 ) );
  BUF_X1 u2_uk_U34 (.Z( u2_uk_n164 ) , .A( u2_uk_n208 ) );
  INV_X1 u2_uk_U350 (.ZN( u2_K10_40 ) , .A( u2_uk_n306 ) );
  AOI22_X1 u2_uk_U351 (.A2( u2_uk_K_r8_2 ) , .B2( u2_uk_K_r8_22 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n306 ) );
  OAI21_X1 u2_uk_U364 (.ZN( u2_K2_33 ) , .A( u2_uk_n1000 ) , .B2( u2_uk_n1258 ) , .B1( u2_uk_n208 ) );
  NAND2_X1 u2_uk_U365 (.A1( u2_uk_K_r0_31 ) , .ZN( u2_uk_n1000 ) , .A2( u2_uk_n147 ) );
  BUF_X1 u2_uk_U37 (.Z( u2_uk_n213 ) , .A( u2_uk_n231 ) );
  BUF_X1 u2_uk_U38 (.Z( u2_uk_n208 ) , .A( u2_uk_n231 ) );
  BUF_X1 u2_uk_U39 (.Z( u2_uk_n214 ) , .A( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U399 (.ZN( u2_K8_16 ) , .B2( u2_uk_n1506 ) , .A2( u2_uk_n1514 ) , .A1( u2_uk_n213 ) , .B1( u2_uk_n27 ) );
  BUF_X1 u2_uk_U40 (.Z( u2_uk_n209 ) , .A( u2_uk_n231 ) );
  OAI22_X1 u2_uk_U412 (.ZN( u2_K12_9 ) , .A1( u2_uk_n100 ) , .B2( u2_uk_n1715 ) , .A2( u2_uk_n1722 ) , .B1( u2_uk_n222 ) );
  INV_X1 u2_uk_U416 (.ZN( u2_K10_37 ) , .A( u2_uk_n299 ) );
  BUF_X1 u2_uk_U42 (.A( u2_uk_n182 ) , .Z( u2_uk_n202 ) );
  BUF_X1 u2_uk_U44 (.A( u2_uk_n182 ) , .Z( u2_uk_n220 ) );
  INV_X1 u2_uk_U446 (.ZN( u2_K10_33 ) , .A( u2_uk_n294 ) );
  AOI22_X1 u2_uk_U447 (.B2( u2_uk_K_r8_22 ) , .A2( u2_uk_K_r8_42 ) , .A1( u2_uk_n117 ) , .B1( u2_uk_n217 ) , .ZN( u2_uk_n294 ) );
  INV_X1 u2_uk_U448 (.ZN( u2_K1_33 ) , .A( u2_uk_n981 ) );
  AOI22_X1 u2_uk_U449 (.B2( u2_key_r_44 ) , .A2( u2_key_r_51 ) , .B1( u2_uk_n100 ) , .A1( u2_uk_n163 ) , .ZN( u2_uk_n981 ) );
  BUF_X1 u2_uk_U46 (.A( u2_uk_n155 ) , .Z( u2_uk_n217 ) );
  OAI22_X1 u2_uk_U472 (.ZN( u2_K1_29 ) , .B2( u2_uk_n1152 ) , .A2( u2_uk_n1158 ) , .B1( u2_uk_n182 ) , .A1( u2_uk_n94 ) );
  BUF_X1 u2_uk_U49 (.Z( u2_uk_n231 ) , .A( u2_uk_n238 ) );
  OAI22_X1 u2_uk_U494 (.ZN( u2_K5_29 ) , .B2( u2_uk_n1377 ) , .A2( u2_uk_n1396 ) , .B1( u2_uk_n148 ) , .A1( u2_uk_n92 ) );
  OAI21_X1 u2_uk_U499 (.ZN( u2_K8_2 ) , .B1( u2_uk_n100 ) , .A( u2_uk_n1105 ) , .B2( u2_uk_n1515 ) );
  OAI22_X1 u2_uk_U501 (.ZN( u2_K5_2 ) , .A2( u2_uk_n1367 ) , .B2( u2_uk_n1372 ) , .B1( u2_uk_n191 ) , .A1( u2_uk_n83 ) );
  OAI21_X1 u2_uk_U514 (.ZN( u2_K8_17 ) , .A( u2_uk_n1101 ) , .B2( u2_uk_n1522 ) , .B1( u2_uk_n187 ) );
  NAND2_X1 u2_uk_U515 (.A1( u2_uk_K_r6_26 ) , .ZN( u2_uk_n1101 ) , .A2( u2_uk_n238 ) );
  OAI21_X1 u2_uk_U523 (.ZN( u2_K12_12 ) , .B2( u2_uk_n1689 ) , .B1( u2_uk_n31 ) , .A( u2_uk_n408 ) );
  OAI21_X1 u2_uk_U527 (.ZN( u2_K5_12 ) , .A( u2_uk_n1041 ) , .B2( u2_uk_n1375 ) , .B1( u2_uk_n163 ) );
  NAND2_X1 u2_uk_U528 (.A1( u2_uk_K_r3_11 ) , .ZN( u2_uk_n1041 ) , .A2( u2_uk_n155 ) );
  OAI22_X1 u2_uk_U533 (.ZN( u2_K1_36 ) , .B2( u2_uk_n1158 ) , .A2( u2_uk_n1165 ) , .B1( u2_uk_n222 ) , .A1( u2_uk_n94 ) );
  OAI22_X1 u2_uk_U553 (.ZN( u2_K1_38 ) , .A1( u2_uk_n10 ) , .B2( u2_uk_n1165 ) , .A2( u2_uk_n1171 ) , .B1( u2_uk_n203 ) );
  INV_X1 u2_uk_U566 (.ZN( u2_K10_38 ) , .A( u2_uk_n301 ) );
  AOI22_X1 u2_uk_U567 (.B2( u2_uk_K_r8_28 ) , .A2( u2_uk_K_r8_8 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n203 ) , .ZN( u2_uk_n301 ) );
  INV_X1 u2_uk_U595 (.ZN( u2_K9_22 ) , .A( u2_uk_n1127 ) );
  AOI22_X1 u2_uk_U596 (.B2( u2_uk_K_r7_41 ) , .A2( u2_uk_K_r7_48 ) , .B1( u2_uk_n109 ) , .ZN( u2_uk_n1127 ) , .A1( u2_uk_n213 ) );
  INV_X1 u2_uk_U600 (.ZN( u2_K5_22 ) , .A( u2_uk_n1044 ) );
  INV_X1 u2_uk_U602 (.ZN( u2_K1_22 ) , .A( u2_uk_n974 ) );
  AOI22_X1 u2_uk_U603 (.B2( u2_key_r_25 ) , .A2( u2_key_r_32 ) , .B1( u2_uk_n109 ) , .A1( u2_uk_n191 ) , .ZN( u2_uk_n974 ) );
  INV_X1 u2_uk_U614 (.ZN( u2_K10_35 ) , .A( u2_uk_n297 ) );
  AOI22_X1 u2_uk_U615 (.B2( u2_uk_K_r8_2 ) , .A2( u2_uk_K_r8_37 ) , .B1( u2_uk_n117 ) , .A1( u2_uk_n238 ) , .ZN( u2_uk_n297 ) );
  INV_X1 u2_uk_U621 (.ZN( u2_K1_35 ) , .A( u2_uk_n982 ) );
  AOI22_X1 u2_uk_U622 (.B2( u2_key_r_28 ) , .A2( u2_key_r_35 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n207 ) , .ZN( u2_uk_n982 ) );
  INV_X1 u2_uk_U644 (.ZN( u2_K1_44 ) , .A( u2_uk_n987 ) );
  AOI22_X1 u2_uk_U645 (.B2( u2_key_r_36 ) , .A2( u2_key_r_43 ) , .B1( u2_uk_n102 ) , .A1( u2_uk_n182 ) , .ZN( u2_uk_n987 ) );
  OAI21_X1 u2_uk_U646 (.ZN( u2_K12_6 ) , .B1( u2_uk_n162 ) , .B2( u2_uk_n1702 ) , .A( u2_uk_n518 ) );
  NAND2_X1 u2_uk_U647 (.A1( u2_uk_K_r10_10 ) , .A2( u2_uk_n148 ) , .ZN( u2_uk_n518 ) );
  INV_X1 u2_uk_U650 (.A( u2_key_r_44 ) , .ZN( u2_uk_n1178 ) );
  OAI22_X1 u2_uk_U651 (.ZN( u2_K14_43 ) , .B1( u2_uk_n142 ) , .B2( u2_uk_n1799 ) , .A2( u2_uk_n1802 ) , .A1( u2_uk_n99 ) );
  OAI21_X1 u2_uk_U665 (.ZN( u2_K14_45 ) , .B2( u2_uk_n1800 ) , .B1( u2_uk_n238 ) , .A( u2_uk_n930 ) );
  NAND2_X1 u2_uk_U666 (.A1( u2_uk_K_r12_16 ) , .A2( u2_uk_n220 ) , .ZN( u2_uk_n930 ) );
  OAI21_X1 u2_uk_U699 (.ZN( u2_K5_7 ) , .A( u2_uk_n1057 ) , .B2( u2_uk_n1405 ) , .B1( u2_uk_n214 ) );
  NAND2_X1 u2_uk_U700 (.A1( u2_uk_K_r3_19 ) , .ZN( u2_uk_n1057 ) , .A2( u2_uk_n217 ) );
  INV_X1 u2_uk_U703 (.ZN( u2_K1_25 ) , .A( u2_uk_n975 ) );
  AOI22_X1 u2_uk_U704 (.B2( u2_key_r_29 ) , .A2( u2_key_r_36 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n975 ) );
  OAI22_X1 u2_uk_U736 (.ZN( u2_K2_42 ) , .B2( u2_uk_n1266 ) , .A2( u2_uk_n1274 ) , .A1( u2_uk_n209 ) , .B1( u2_uk_n60 ) );
  INV_X1 u2_uk_U739 (.ZN( u2_K1_42 ) , .A( u2_uk_n986 ) );
  OAI22_X1 u2_uk_U750 (.ZN( u2_K8_13 ) , .A2( u2_uk_n1501 ) , .B2( u2_uk_n1507 ) , .B1( u2_uk_n231 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U761 (.ZN( u2_K9_21 ) , .A1( u2_uk_n117 ) , .B2( u2_uk_n1568 ) , .A2( u2_uk_n1573 ) , .B1( u2_uk_n208 ) );
  INV_X1 u2_uk_U785 (.ZN( u2_K5_27 ) , .A( u2_uk_n1046 ) );
  INV_X1 u2_uk_U791 (.ZN( u2_K1_27 ) , .A( u2_uk_n977 ) );
  AOI22_X1 u2_uk_U792 (.B2( u2_key_r_14 ) , .A2( u2_key_r_21 ) , .B1( u2_uk_n128 ) , .A1( u2_uk_n162 ) , .ZN( u2_uk_n977 ) );
  INV_X1 u2_uk_U793 (.ZN( u2_K9_27 ) , .A( u2_uk_n1129 ) );
  AOI22_X1 u2_uk_U794 (.B2( u2_uk_K_r7_2 ) , .A2( u2_uk_K_r7_9 ) , .B1( u2_uk_n109 ) , .ZN( u2_uk_n1129 ) , .A1( u2_uk_n163 ) );
  OAI22_X1 u2_uk_U828 (.ZN( u2_K8_6 ) , .B2( u2_uk_n1514 ) , .A2( u2_uk_n1519 ) , .A1( u2_uk_n188 ) , .B1( u2_uk_n83 ) );
  INV_X1 u2_uk_U831 (.ZN( u2_K12_3 ) , .A( u2_uk_n500 ) );
  OAI22_X1 u2_uk_U844 (.ZN( u2_K1_1 ) , .A1( u2_uk_n11 ) , .B2( u2_uk_n1174 ) , .A2( u2_uk_n1179 ) , .B1( u2_uk_n182 ) );
  OAI22_X1 u2_uk_U859 (.ZN( u2_K12_10 ) , .B1( u2_uk_n10 ) , .B2( u2_uk_n1688 ) , .A2( u2_uk_n1709 ) , .A1( u2_uk_n207 ) );
  INV_X1 u2_uk_U86 (.ZN( u2_K2_41 ) , .A( u2_uk_n1001 ) );
  OAI22_X1 u2_uk_U860 (.ZN( u2_K12_11 ) , .A1( u2_uk_n146 ) , .A2( u2_uk_n1683 ) , .B2( u2_uk_n1709 ) , .B1( u2_uk_n63 ) );
  OAI22_X1 u2_uk_U870 (.ZN( u2_K8_1 ) , .A2( u2_uk_n1502 ) , .B2( u2_uk_n1518 ) , .A1( u2_uk_n182 ) , .B1( u2_uk_n27 ) );
  OAI22_X1 u2_uk_U881 (.ZN( u2_K9_24 ) , .B1( u2_uk_n128 ) , .B2( u2_uk_n1544 ) , .A2( u2_uk_n1586 ) , .A1( u2_uk_n220 ) );
  OAI22_X1 u2_uk_U905 (.ZN( u2_K2_39 ) , .B1( u2_uk_n11 ) , .A2( u2_uk_n1236 ) , .B2( u2_uk_n1251 ) , .A1( u2_uk_n164 ) );
  OAI22_X1 u2_uk_U924 (.ZN( u2_K14_47 ) , .B1( u2_uk_n145 ) , .B2( u2_uk_n1790 ) , .A2( u2_uk_n1800 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U945 (.ZN( u2_K2_38 ) , .B2( u2_uk_n1246 ) , .A2( u2_uk_n1265 ) , .B1( u2_uk_n129 ) , .A1( u2_uk_n92 ) );
  OAI22_X1 u2_uk_U947 (.ZN( u2_K2_37 ) , .A2( u2_uk_n1237 ) , .B2( u2_uk_n1264 ) , .B1( u2_uk_n129 ) , .A1( u2_uk_n93 ) );
  OAI22_X1 u2_uk_U965 (.ZN( u2_K1_34 ) , .A1( u2_uk_n100 ) , .B2( u2_uk_n1144 ) , .A2( u2_uk_n1149 ) , .B1( u2_uk_n147 ) );
  OAI22_X1 u2_uk_U966 (.ZN( u2_K1_47 ) , .B2( u2_uk_n1142 ) , .A2( u2_uk_n1147 ) , .B1( u2_uk_n142 ) , .A1( u2_uk_n99 ) );
  OAI22_X1 u2_uk_U98 (.ZN( u2_K12_5 ) , .A2( u2_uk_n1682 ) , .B2( u2_uk_n1708 ) , .A1( u2_uk_n202 ) , .B1( u2_uk_n94 ) );
  OAI21_X1 u2_uk_U983 (.ZN( u2_K14_46 ) , .B1( u2_uk_n102 ) , .B2( u2_uk_n1790 ) , .A( u2_uk_n931 ) );
  OAI21_X1 u2_uk_U989 (.ZN( u2_K8_4 ) , .B1( u2_uk_n102 ) , .A( u2_uk_n1116 ) , .B2( u2_uk_n1507 ) );
  OAI21_X1 u2_uk_U991 (.ZN( u2_K5_4 ) , .A( u2_uk_n1055 ) , .B1( u2_uk_n110 ) , .B2( u2_uk_n1381 ) );
  NAND2_X1 u2_uk_U992 (.A1( u2_uk_K_r3_4 ) , .ZN( u2_uk_n1055 ) , .A2( u2_uk_n63 ) );
endmodule

