module aes_aes_die_4 ( sa03_4, sa03_5, us03_n445, us03_n450, us03_n458, us03_n462, us03_n463, us03_n695, us03_n722, 
       us03_n726, us03_n727, us03_n728, us03_n742, us03_n745, us03_n748, us03_n760, us03_n761, us03_n777, 
       us03_n783, us03_n784, us03_n786, us03_n788, us03_n790, us03_n801, us03_n803, us03_n804, us03_n811, 
       us03_n812, us03_n813, us03_n814, us03_n815, sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7 );
  input sa03_4, sa03_5, us03_n445, us03_n450, us03_n458, us03_n462, us03_n463, us03_n695, us03_n722, 
        us03_n726, us03_n727, us03_n728, us03_n742, us03_n745, us03_n748, us03_n760, us03_n761, us03_n777, 
        us03_n783, us03_n784, us03_n786, us03_n788, us03_n790, us03_n801, us03_n803, us03_n804, us03_n811, 
        us03_n812, us03_n813, us03_n814, us03_n815;
  output sa03_sr_0, sa03_sr_1, sa03_sr_2, sa03_sr_3, sa03_sr_4, sa03_sr_5, sa03_sr_6, sa03_sr_7;
  wire us03_n438, us03_n439, us03_n440, us03_n441, us03_n442, us03_n443, us03_n444, us03_n448, us03_n454, 
       us03_n455, us03_n456, us03_n457, us03_n461, us03_n464, us03_n465, us03_n466, us03_n467, us03_n468, 
       us03_n471, us03_n472, us03_n473, us03_n474, us03_n475, us03_n476, us03_n477, us03_n478, us03_n479, 
       us03_n480, us03_n481, us03_n482, us03_n483, us03_n484, us03_n485, us03_n486, us03_n487, us03_n488, 
       us03_n489, us03_n490, us03_n491, us03_n492, us03_n493, us03_n494, us03_n495, us03_n496, us03_n497, 
       us03_n498, us03_n499, us03_n500, us03_n501, us03_n502, us03_n503, us03_n504, us03_n505, us03_n506, 
       us03_n507, us03_n508, us03_n509, us03_n510, us03_n511, us03_n512, us03_n513, us03_n514, us03_n515, 
       us03_n516, us03_n517, us03_n518, us03_n519, us03_n520, us03_n521, us03_n522, us03_n523, us03_n524, 
       us03_n525, us03_n526, us03_n527, us03_n528, us03_n529, us03_n530, us03_n531, us03_n532, us03_n533, 
       us03_n534, us03_n535, us03_n536, us03_n537, us03_n538, us03_n539, us03_n540, us03_n541, us03_n542, 
       us03_n543, us03_n544, us03_n545, us03_n546, us03_n547, us03_n548, us03_n549, us03_n550, us03_n551, 
       us03_n552, us03_n553, us03_n554, us03_n555, us03_n556, us03_n557, us03_n558, us03_n559, us03_n560, 
       us03_n561, us03_n562, us03_n563, us03_n564, us03_n565, us03_n566, us03_n567, us03_n568, us03_n569, 
       us03_n570, us03_n571, us03_n572, us03_n573, us03_n574, us03_n575, us03_n576, us03_n577, us03_n578, 
       us03_n579, us03_n580, us03_n581, us03_n582, us03_n583, us03_n584, us03_n585, us03_n586, us03_n587, 
       us03_n588, us03_n589, us03_n590, us03_n591, us03_n592, us03_n593, us03_n594, us03_n595, us03_n596, 
       us03_n597, us03_n598, us03_n599, us03_n600, us03_n601, us03_n602, us03_n603, us03_n604, us03_n605, 
       us03_n606, us03_n607, us03_n608, us03_n609, us03_n610, us03_n611, us03_n612, us03_n613, us03_n614, 
       us03_n615, us03_n616, us03_n617, us03_n618, us03_n619, us03_n620, us03_n621, us03_n622, us03_n623, 
       us03_n624, us03_n625, us03_n626, us03_n627, us03_n628, us03_n629, us03_n630, us03_n631, us03_n632, 
       us03_n633, us03_n634, us03_n635, us03_n636, us03_n637, us03_n638, us03_n639, us03_n640, us03_n641, 
       us03_n642, us03_n643, us03_n644, us03_n645, us03_n646, us03_n647, us03_n648, us03_n649, us03_n650, 
       us03_n651, us03_n652, us03_n653, us03_n654, us03_n655, us03_n656, us03_n657, us03_n658, us03_n659, 
       us03_n660, us03_n661, us03_n662, us03_n663, us03_n664, us03_n665, us03_n666, us03_n667, us03_n668, 
       us03_n669, us03_n670, us03_n671, us03_n672, us03_n673, us03_n674, us03_n675, us03_n676, us03_n677, 
       us03_n678, us03_n679, us03_n680, us03_n681, us03_n682, us03_n683, us03_n684, us03_n685, us03_n686, 
       us03_n687, us03_n688, us03_n689, us03_n690, us03_n691, us03_n692, us03_n693, us03_n694, us03_n696, 
       us03_n697, us03_n698, us03_n699, us03_n700, us03_n701, us03_n702, us03_n703, us03_n704, us03_n705, 
       us03_n706, us03_n707, us03_n708, us03_n709, us03_n710, us03_n711, us03_n712, us03_n713, us03_n714, 
       us03_n715, us03_n716, us03_n717, us03_n718, us03_n719, us03_n720, us03_n721, us03_n723, us03_n724, 
       us03_n725, us03_n729, us03_n730, us03_n731, us03_n732, us03_n733, us03_n734, us03_n735, us03_n736, 
       us03_n737, us03_n738, us03_n739, us03_n740, us03_n741, us03_n743, us03_n744, us03_n746, us03_n747, 
       us03_n749, us03_n750, us03_n751, us03_n752, us03_n753, us03_n754, us03_n755, us03_n756, us03_n757, 
       us03_n758, us03_n759, us03_n762, us03_n763, us03_n764, us03_n765, us03_n766, us03_n767, us03_n768, 
       us03_n769, us03_n770, us03_n771, us03_n772, us03_n773, us03_n774, us03_n775, us03_n776, us03_n778, 
       us03_n779, us03_n780, us03_n781, us03_n782, us03_n785, us03_n787, us03_n789, us03_n791, us03_n792, 
       us03_n793, us03_n794, us03_n795, us03_n796, us03_n797, us03_n798, us03_n799, us03_n800, us03_n802, 
       us03_n805, us03_n806, us03_n807, us03_n808, us03_n809, us03_n810, us03_n816, us03_n817, us03_n818, 
       us03_n819, us03_n820, us03_n821, us03_n822, us03_n823, us03_n828, us03_n829, us03_n830, us03_n831, 
       us03_n832, us03_n833, us03_n834, us03_n835, us03_n836, us03_n837, us03_n838, us03_n839, us03_n840, 
       us03_n841, us03_n842, us03_n843, us03_n844, us03_n848, us03_n849, us03_n850, us03_n851, us03_n852, 
       us03_n853, us03_n854, us03_n855, us03_n857, us03_n858, us03_n859, us03_n860, us03_n861, us03_n862, 
       us03_n863, us03_n864, us03_n865, us03_n866, us03_n867, us03_n868, us03_n869, us03_n870, us03_n871, 
       us03_n872, us03_n873,  us03_n874;
  INV_X1 us03_U10 (.A( us03_n678 ) , .ZN( us03_n838 ) );
  NOR4_X1 us03_U100 (.A4( us03_n607 ) , .A3( us03_n608 ) , .A2( us03_n609 ) , .A1( us03_n610 ) , .ZN( us03_n617 ) );
  NOR4_X1 us03_U101 (.A4( us03_n612 ) , .A3( us03_n613 ) , .A2( us03_n614 ) , .A1( us03_n615 ) , .ZN( us03_n616 ) );
  NOR2_X1 us03_U102 (.ZN( us03_n684 ) , .A1( us03_n829 ) , .A2( us03_n830 ) );
  NAND4_X1 us03_U103 (.A4( us03_n471 ) , .A3( us03_n472 ) , .A2( us03_n473 ) , .A1( us03_n474 ) , .ZN( us03_n676 ) );
  NOR4_X1 us03_U104 (.A4( us03_n468 ) , .ZN( us03_n474 ) , .A3( us03_n554 ) , .A1( us03_n733 ) , .A2( us03_n753 ) );
  NOR4_X1 us03_U105 (.ZN( us03_n473 ) , .A1( us03_n529 ) , .A3( us03_n566 ) , .A4( us03_n598 ) , .A2( us03_n640 ) );
  NOR4_X1 us03_U106 (.ZN( us03_n472 ) , .A1( us03_n504 ) , .A3( us03_n542 ) , .A2( us03_n581 ) , .A4( us03_n714 ) );
  NAND4_X1 us03_U107 (.ZN( sa03_sr_1 ) , .A4( us03_n593 ) , .A3( us03_n594 ) , .A2( us03_n595 ) , .A1( us03_n596 ) );
  AOI211_X1 us03_U108 (.B( us03_n587 ) , .A( us03_n588 ) , .ZN( us03_n594 ) , .C2( us03_n809 ) , .C1( us03_n831 ) );
  NOR4_X1 us03_U109 (.A4( us03_n589 ) , .A3( us03_n590 ) , .A2( us03_n591 ) , .A1( us03_n592 ) , .ZN( us03_n593 ) );
  NOR4_X1 us03_U11 (.A4( us03_n443 ) , .A3( us03_n444 ) , .A2( us03_n514 ) , .A1( us03_n539 ) , .ZN( us03_n704 ) );
  AOI211_X1 us03_U110 (.A( us03_n586 ) , .ZN( us03_n595 ) , .B( us03_n619 ) , .C1( us03_n843 ) , .C2( us03_n853 ) );
  NAND4_X1 us03_U111 (.ZN( sa03_sr_0 ) , .A4( us03_n499 ) , .A3( us03_n500 ) , .A2( us03_n501 ) , .A1( us03_n502 ) );
  NOR4_X1 us03_U112 (.A4( us03_n496 ) , .A3( us03_n497 ) , .A2( us03_n498 ) , .ZN( us03_n499 ) , .A1( us03_n525 ) );
  AOI221_X1 us03_U113 (.A( us03_n495 ) , .ZN( us03_n500 ) , .B2( us03_n841 ) , .C1( us03_n844 ) , .C2( us03_n858 ) , .B1( us03_n860 ) );
  AOI211_X1 us03_U114 (.A( us03_n494 ) , .ZN( us03_n501 ) , .B( us03_n800 ) , .C2( us03_n837 ) , .C1( us03_n849 ) );
  NAND4_X1 us03_U115 (.A4( us03_n689 ) , .A3( us03_n690 ) , .A1( us03_n691 ) , .ZN( us03_n774 ) , .A2( us03_n870 ) );
  INV_X1 us03_U116 (.A( us03_n677 ) , .ZN( us03_n870 ) );
  AOI221_X1 us03_U117 (.A( us03_n679 ) , .ZN( us03_n690 ) , .B2( us03_n838 ) , .C1( us03_n840 ) , .C2( us03_n860 ) , .B1( us03_n863 ) );
  NOR4_X1 us03_U118 (.A4( us03_n685 ) , .A3( us03_n686 ) , .A2( us03_n687 ) , .A1( us03_n688 ) , .ZN( us03_n689 ) );
  NOR2_X1 us03_U119 (.ZN( us03_n731 ) , .A2( us03_n830 ) , .A1( us03_n843 ) );
  OR3_X1 us03_U12 (.ZN( us03_n444 ) , .A1( us03_n526 ) , .A3( us03_n575 ) , .A2( us03_n873 ) );
  NAND4_X1 us03_U120 (.A4( us03_n717 ) , .A3( us03_n718 ) , .A2( us03_n719 ) , .ZN( us03_n739 ) , .A1( us03_n855 ) );
  INV_X1 us03_U121 (.A( us03_n707 ) , .ZN( us03_n855 ) );
  NOR4_X1 us03_U122 (.A4( us03_n713 ) , .A3( us03_n714 ) , .A2( us03_n715 ) , .A1( us03_n716 ) , .ZN( us03_n717 ) );
  AOI221_X1 us03_U123 (.A( us03_n708 ) , .ZN( us03_n719 ) , .C2( us03_n842 ) , .B2( us03_n843 ) , .C1( us03_n859 ) , .B1( us03_n860 ) );
  NOR2_X1 us03_U124 (.ZN( us03_n645 ) , .A1( us03_n852 ) , .A2( us03_n866 ) );
  NAND4_X1 us03_U125 (.A4( us03_n571 ) , .A3( us03_n572 ) , .A1( us03_n573 ) , .ZN( us03_n721 ) , .A2( us03_n872 ) );
  NOR4_X1 us03_U126 (.A4( us03_n567 ) , .A3( us03_n568 ) , .A2( us03_n569 ) , .A1( us03_n570 ) , .ZN( us03_n571 ) );
  AOI221_X1 us03_U127 (.A( us03_n562 ) , .C2( us03_n563 ) , .ZN( us03_n572 ) , .B2( us03_n843 ) , .B1( us03_n850 ) , .C1( us03_n851 ) );
  INV_X1 us03_U128 (.A( us03_n605 ) , .ZN( us03_n872 ) );
  NAND4_X1 us03_U129 (.A4( us03_n491 ) , .A3( us03_n492 ) , .A1( us03_n493 ) , .ZN( us03_n800 ) , .A2( us03_n865 ) );
  OR4_X1 us03_U13 (.A4( us03_n440 ) , .A2( us03_n441 ) , .A1( us03_n442 ) , .ZN( us03_n443 ) , .A3( us03_n551 ) );
  AOI221_X1 us03_U130 (.A( us03_n487 ) , .ZN( us03_n492 ) , .B2( us03_n834 ) , .C2( us03_n839 ) , .C1( us03_n849 ) , .B1( us03_n858 ) );
  INV_X1 us03_U131 (.A( us03_n776 ) , .ZN( us03_n865 ) );
  NOR2_X1 us03_U132 (.ZN( us03_n493 ) , .A1( us03_n676 ) , .A2( us03_n692 ) );
  INV_X1 us03_U133 (.A( us03_n760 ) , .ZN( us03_n828 ) );
  INV_X1 us03_U134 (.A( us03_n461 ) , .ZN( us03_n862 ) );
  OAI21_X1 us03_U135 (.ZN( us03_n461 ) , .B1( us03_n807 ) , .A( us03_n832 ) , .B2( us03_n849 ) );
  OR4_X1 us03_U136 (.A4( us03_n578 ) , .A3( us03_n579 ) , .A2( us03_n580 ) , .A1( us03_n581 ) , .ZN( us03_n582 ) );
  OR4_X1 us03_U137 (.A4( us03_n564 ) , .A3( us03_n565 ) , .A2( us03_n566 ) , .ZN( us03_n570 ) , .A1( us03_n663 ) );
  OR4_X1 us03_U138 (.A4( us03_n516 ) , .A2( us03_n517 ) , .A1( us03_n518 ) , .ZN( us03_n520 ) , .A3( us03_n819 ) );
  OR4_X1 us03_U139 (.A4( us03_n680 ) , .A3( us03_n681 ) , .A2( us03_n682 ) , .A1( us03_n683 ) , .ZN( us03_n688 ) );
  INV_X1 us03_U14 (.A( us03_n611 ) , .ZN( us03_n873 ) );
  OR4_X1 us03_U140 (.ZN( us03_n464 ) , .A4( us03_n516 ) , .A3( us03_n527 ) , .A2( us03_n576 ) , .A1( us03_n710 ) );
  NAND2_X1 us03_U141 (.ZN( us03_n611 ) , .A2( us03_n835 ) , .A1( us03_n871 ) );
  OR3_X1 us03_U142 (.A3( us03_n504 ) , .A2( us03_n505 ) , .A1( us03_n506 ) , .ZN( us03_n509 ) );
  AOI221_X1 us03_U143 (.A( us03_n711 ) , .B2( us03_n712 ) , .ZN( us03_n718 ) , .C1( us03_n830 ) , .B1( us03_n837 ) , .C2( us03_n861 ) );
  OR2_X1 us03_U144 (.A2( us03_n709 ) , .A1( us03_n710 ) , .ZN( us03_n711 ) );
  INV_X1 us03_U145 (.A( us03_n752 ) , .ZN( us03_n867 ) );
  OAI21_X1 us03_U146 (.B1( us03_n751 ) , .ZN( us03_n752 ) , .A( us03_n843 ) , .B2( us03_n866 ) );
  INV_X1 us03_U147 (.A( us03_n670 ) , .ZN( us03_n857 ) );
  AOI21_X1 us03_U148 (.A( us03_n668 ) , .B1( us03_n669 ) , .ZN( us03_n670 ) , .B2( us03_n854 ) );
  AOI222_X1 us03_U149 (.ZN( us03_n658 ) , .A2( us03_n837 ) , .B1( us03_n839 ) , .C2( us03_n843 ) , .A1( us03_n858 ) , .C1( us03_n861 ) , .B2( us03_n868 ) );
  INV_X1 us03_U15 (.A( us03_n747 ) , .ZN( us03_n861 ) );
  INV_X1 us03_U150 (.A( us03_n645 ) , .ZN( us03_n868 ) );
  OAI22_X1 us03_U151 (.ZN( us03_n481 ) , .A1( us03_n706 ) , .B2( us03_n783 ) , .A2( us03_n804 ) , .B1( us03_n810 ) );
  NAND2_X1 us03_U152 (.A1( us03_n445 ) , .A2( us03_n463 ) , .ZN( us03_n747 ) );
  OAI222_X1 us03_U153 (.B2( us03_n745 ) , .B1( us03_n746 ) , .A2( us03_n747 ) , .ZN( us03_n755 ) , .C2( us03_n803 ) , .C1( us03_n812 ) , .A1( us03_n815 ) );
  OAI222_X1 us03_U154 (.B2( us03_n706 ) , .ZN( us03_n707 ) , .C2( us03_n722 ) , .B1( us03_n745 ) , .A1( us03_n804 ) , .C1( us03_n812 ) , .A2( us03_n813 ) );
  OAI222_X1 us03_U155 (.ZN( us03_n615 ) , .B1( us03_n695 ) , .C1( us03_n722 ) , .C2( us03_n745 ) , .B2( us03_n784 ) , .A2( us03_n790 ) , .A1( us03_n814 ) );
  OAI222_X1 us03_U156 (.ZN( us03_n503 ) , .C2( us03_n623 ) , .B2( us03_n645 ) , .B1( us03_n745 ) , .A2( us03_n746 ) , .C1( us03_n803 ) , .A1( us03_n804 ) );
  AOI22_X1 us03_U157 (.ZN( us03_n694 ) , .A1( us03_n828 ) , .B2( us03_n841 ) , .A2( us03_n863 ) , .B1( us03_n866 ) );
  INV_X1 us03_U158 (.A( us03_n728 ) , .ZN( us03_n837 ) );
  AOI221_X1 us03_U159 (.A( us03_n762 ) , .ZN( us03_n772 ) , .C2( us03_n808 ) , .B2( us03_n833 ) , .C1( us03_n853 ) , .B1( us03_n864 ) );
  AOI222_X1 us03_U16 (.ZN( us03_n561 ) , .B1( us03_n828 ) , .C1( us03_n839 ) , .A2( us03_n841 ) , .A1( us03_n852 ) , .B2( us03_n861 ) , .C2( us03_n871 ) );
  AOI21_X1 us03_U160 (.B2( us03_n761 ) , .ZN( us03_n762 ) , .A( us03_n786 ) , .B1( us03_n790 ) );
  INV_X1 us03_U161 (.A( us03_n759 ) , .ZN( us03_n833 ) );
  INV_X1 us03_U163 (.A( us03_n788 ) , .ZN( us03_n830 ) );
  OAI22_X1 us03_U164 (.ZN( us03_n635 ) , .A1( us03_n697 ) , .B2( us03_n726 ) , .A2( us03_n760 ) , .B1( us03_n814 ) );
  OAI221_X1 us03_U165 (.A( us03_n725 ) , .C2( us03_n726 ) , .B2( us03_n727 ) , .B1( us03_n728 ) , .ZN( us03_n735 ) , .C1( us03_n815 ) );
  AOI22_X1 us03_U166 (.ZN( us03_n725 ) , .B1( us03_n830 ) , .A2( us03_n836 ) , .A1( us03_n861 ) , .B2( us03_n864 ) );
  OAI22_X1 us03_U167 (.ZN( us03_n487 ) , .A1( us03_n722 ) , .B2( us03_n726 ) , .B1( us03_n728 ) , .A2( us03_n777 ) );
  OAI22_X1 us03_U168 (.ZN( us03_n622 ) , .B1( us03_n667 ) , .B2( us03_n745 ) , .A1( us03_n813 ) , .A2( us03_n814 ) );
  OAI22_X1 us03_U169 (.A1( us03_n722 ) , .ZN( us03_n724 ) , .B2( us03_n748 ) , .B1( us03_n810 ) , .A2( us03_n814 ) );
  NOR4_X1 us03_U17 (.ZN( us03_n471 ) , .A2( us03_n519 ) , .A4( us03_n592 ) , .A1( us03_n607 ) , .A3( us03_n627 ) );
  OAI22_X1 us03_U170 (.B2( us03_n777 ) , .B1( us03_n778 ) , .ZN( us03_n779 ) , .A2( us03_n812 ) , .A1( us03_n813 ) );
  OAI22_X1 us03_U171 (.B2( us03_n742 ) , .ZN( us03_n744 ) , .A2( us03_n760 ) , .B1( us03_n778 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U172 (.B2( us03_n801 ) , .B1( us03_n802 ) , .A2( us03_n803 ) , .A1( us03_n804 ) , .ZN( us03_n806 ) );
  OAI22_X1 us03_U173 (.ZN( us03_n494 ) , .A2( us03_n742 ) , .A1( us03_n778 ) , .B1( us03_n789 ) , .B2( us03_n804 ) );
  INV_X1 us03_U174 (.A( us03_n742 ) , .ZN( us03_n835 ) );
  INV_X1 us03_U175 (.A( us03_n814 ) , .ZN( us03_n829 ) );
  INV_X1 us03_U176 (.A( us03_n786 ) , .ZN( us03_n843 ) );
  INV_X1 us03_U177 (.A( us03_n812 ) , .ZN( us03_n831 ) );
  OAI22_X1 us03_U178 (.ZN( us03_n588 ) , .B1( us03_n728 ) , .B2( us03_n747 ) , .A2( us03_n784 ) , .A1( us03_n801 ) );
  OAI22_X1 us03_U179 (.ZN( us03_n693 ) , .A2( us03_n728 ) , .A1( us03_n778 ) , .B1( us03_n789 ) , .B2( us03_n815 ) );
  NOR4_X1 us03_U18 (.ZN( us03_n477 ) , .A1( us03_n518 ) , .A4( us03_n555 ) , .A3( us03_n580 ) , .A2( us03_n628 ) );
  OAI22_X1 us03_U180 (.ZN( us03_n708 ) , .A2( us03_n726 ) , .B2( us03_n727 ) , .A1( us03_n742 ) , .B1( us03_n811 ) );
  INV_X1 us03_U181 (.A( us03_n667 ) , .ZN( us03_n863 ) );
  NOR2_X1 us03_U182 (.A1( us03_n695 ) , .ZN( us03_n768 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U183 (.ZN( us03_n664 ) , .A1( us03_n726 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U184 (.ZN( us03_n592 ) , .A2( us03_n695 ) , .A1( us03_n726 ) );
  NOR2_X1 us03_U185 (.ZN( us03_n568 ) , .A1( us03_n726 ) , .A2( us03_n804 ) );
  NOR2_X1 us03_U186 (.ZN( us03_n716 ) , .A2( us03_n722 ) , .A1( us03_n742 ) );
  NOR2_X1 us03_U187 (.ZN( us03_n544 ) , .A2( us03_n778 ) , .A1( us03_n812 ) );
  NOR2_X1 us03_U188 (.ZN( us03_n575 ) , .A2( us03_n697 ) , .A1( us03_n812 ) );
  NOR2_X1 us03_U189 (.ZN( us03_n652 ) , .A1( us03_n726 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U19 (.A4( us03_n530 ) , .A3( us03_n531 ) , .A2( us03_n532 ) , .ZN( us03_n533 ) , .A1( us03_n818 ) );
  NOR2_X1 us03_U190 (.ZN( us03_n610 ) , .A1( us03_n777 ) , .A2( us03_n784 ) );
  INV_X1 us03_U191 (.A( us03_n748 ) , .ZN( us03_n840 ) );
  NOR2_X1 us03_U192 (.ZN( us03_n530 ) , .A2( us03_n747 ) , .A1( us03_n748 ) );
  NOR2_X1 us03_U193 (.ZN( us03_n627 ) , .A2( us03_n726 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U194 (.ZN( us03_n613 ) , .A1( us03_n783 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U195 (.ZN( us03_n599 ) , .A2( us03_n778 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U196 (.ZN( us03_n609 ) , .A2( us03_n778 ) , .A1( us03_n804 ) );
  INV_X1 us03_U197 (.A( us03_n745 ) , .ZN( us03_n832 ) );
  NOR2_X1 us03_U198 (.A2( us03_n742 ) , .ZN( us03_n767 ) , .A1( us03_n810 ) );
  NOR2_X1 us03_U199 (.ZN( us03_n526 ) , .A2( us03_n722 ) , .A1( us03_n801 ) );
  NOR4_X1 us03_U20 (.ZN( us03_n454 ) , .A2( us03_n515 ) , .A1( us03_n541 ) , .A3( us03_n577 ) , .A4( us03_n613 ) );
  NOR2_X1 us03_U200 (.ZN( us03_n529 ) , .A2( us03_n778 ) , .A1( us03_n814 ) );
  NOR2_X1 us03_U201 (.ZN( us03_n626 ) , .A2( us03_n667 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U202 (.ZN( us03_n597 ) , .A2( us03_n789 ) , .A1( us03_n814 ) );
  INV_X1 us03_U203 (.A( us03_n790 ) , .ZN( us03_n849 ) );
  NOR2_X1 us03_U204 (.ZN( us03_n650 ) , .A1( us03_n667 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U205 (.A1( us03_n667 ) , .ZN( us03_n671 ) , .A2( us03_n742 ) );
  NOR2_X1 us03_U206 (.ZN( us03_n600 ) , .A1( us03_n667 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U207 (.A1( us03_n667 ) , .ZN( us03_n686 ) , .A2( us03_n814 ) );
  NOR2_X1 us03_U208 (.A2( us03_n706 ) , .A1( us03_n748 ) , .ZN( us03_n769 ) );
  NOR2_X1 us03_U209 (.A1( us03_n667 ) , .ZN( us03_n764 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U21 (.A4( us03_n539 ) , .A3( us03_n540 ) , .A2( us03_n541 ) , .ZN( us03_n548 ) , .A1( us03_n686 ) );
  NOR2_X1 us03_U210 (.A1( us03_n697 ) , .ZN( us03_n766 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U211 (.ZN( us03_n539 ) , .A2( us03_n695 ) , .A1( us03_n697 ) );
  NOR2_X1 us03_U212 (.ZN( us03_n525 ) , .A1( us03_n667 ) , .A2( us03_n777 ) );
  NOR2_X1 us03_U213 (.ZN( us03_n665 ) , .A1( us03_n748 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U214 (.ZN( us03_n553 ) , .A1( us03_n748 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U215 (.ZN( us03_n506 ) , .A2( us03_n778 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U216 (.ZN( us03_n541 ) , .A2( us03_n706 ) , .A1( us03_n783 ) );
  NOR2_X1 us03_U217 (.ZN( us03_n662 ) , .A1( us03_n783 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U218 (.A2( us03_n695 ) , .ZN( us03_n714 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U219 (.B1( us03_n438 ) , .ZN( us03_n442 ) , .A2( us03_n726 ) , .A1( us03_n742 ) , .B2( us03_n747 ) );
  NOR2_X1 us03_U22 (.ZN( us03_n678 ) , .A2( us03_n832 ) , .A1( us03_n837 ) );
  NOR3_X1 us03_U220 (.ZN( us03_n438 ) , .A2( us03_n834 ) , .A3( us03_n835 ) , .A1( us03_n844 ) );
  NOR2_X1 us03_U221 (.ZN( us03_n505 ) , .A1( us03_n810 ) , .A2( us03_n815 ) );
  INV_X1 us03_U222 (.A( us03_n804 ) , .ZN( us03_n839 ) );
  NOR2_X1 us03_U223 (.ZN( us03_n659 ) , .A1( us03_n727 ) , .A2( us03_n788 ) );
  NOR2_X1 us03_U224 (.ZN( us03_n660 ) , .A2( us03_n695 ) , .A1( us03_n727 ) );
  NOR2_X1 us03_U225 (.ZN( us03_n555 ) , .A1( us03_n790 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U226 (.ZN( us03_n543 ) , .A1( us03_n747 ) , .A2( us03_n812 ) );
  NOR2_X1 us03_U227 (.ZN( us03_n507 ) , .A1( us03_n727 ) , .A2( us03_n777 ) );
  INV_X1 us03_U228 (.A( us03_n801 ) , .ZN( us03_n841 ) );
  NOR2_X1 us03_U229 (.A2( us03_n695 ) , .A1( us03_n778 ) , .ZN( us03_n818 ) );
  NOR4_X1 us03_U23 (.A4( us03_n512 ) , .A3( us03_n513 ) , .A2( us03_n514 ) , .A1( us03_n515 ) , .ZN( us03_n522 ) );
  NOR2_X1 us03_U230 (.ZN( us03_n528 ) , .A2( us03_n742 ) , .A1( us03_n790 ) );
  OAI22_X1 us03_U231 (.B2( us03_n748 ) , .B1( us03_n749 ) , .A1( us03_n750 ) , .ZN( us03_n754 ) , .A2( us03_n804 ) );
  NOR2_X1 us03_U232 (.ZN( us03_n749 ) , .A2( us03_n850 ) , .A1( us03_n858 ) );
  NOR3_X1 us03_U233 (.ZN( us03_n750 ) , .A2( us03_n851 ) , .A1( us03_n861 ) , .A3( us03_n863 ) );
  NOR2_X1 us03_U234 (.A1( us03_n747 ) , .ZN( us03_n765 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U235 (.A2( us03_n742 ) , .ZN( us03_n753 ) , .A1( us03_n803 ) );
  NOR2_X1 us03_U236 (.ZN( us03_n542 ) , .A2( us03_n783 ) , .A1( us03_n790 ) );
  NOR2_X1 us03_U237 (.ZN( us03_n661 ) , .A1( us03_n727 ) , .A2( us03_n783 ) );
  INV_X1 us03_U238 (.A( us03_n726 ) , .ZN( us03_n850 ) );
  NOR2_X1 us03_U239 (.ZN( us03_n629 ) , .A1( us03_n722 ) , .A2( us03_n811 ) );
  AOI222_X1 us03_U24 (.ZN( us03_n523 ) , .A1( us03_n832 ) , .B2( us03_n835 ) , .C1( us03_n842 ) , .C2( us03_n848 ) , .A2( us03_n850 ) , .B1( us03_n864 ) );
  NOR2_X1 us03_U240 (.ZN( us03_n733 ) , .A2( us03_n801 ) , .A1( us03_n803 ) );
  NOR2_X1 us03_U241 (.ZN( us03_n612 ) , .A1( us03_n760 ) , .A2( us03_n810 ) );
  NOR4_X1 us03_U242 (.A2( us03_n489 ) , .A1( us03_n490 ) , .ZN( us03_n491 ) , .A3( us03_n578 ) , .A4( us03_n610 ) );
  OR4_X1 us03_U243 (.ZN( us03_n490 ) , .A4( us03_n532 ) , .A2( us03_n545 ) , .A1( us03_n557 ) , .A3( us03_n630 ) );
  OAI22_X1 us03_U244 (.B1( us03_n488 ) , .ZN( us03_n489 ) , .A1( us03_n684 ) , .A2( us03_n761 ) , .B2( us03_n815 ) );
  NOR3_X1 us03_U245 (.ZN( us03_n488 ) , .A1( us03_n780 ) , .A2( us03_n848 ) , .A3( us03_n861 ) );
  NOR2_X1 us03_U246 (.ZN( us03_n504 ) , .A2( us03_n726 ) , .A1( us03_n760 ) );
  NOR2_X1 us03_U247 (.ZN( us03_n514 ) , .A1( us03_n706 ) , .A2( us03_n742 ) );
  NOR2_X1 us03_U248 (.ZN( us03_n715 ) , .A2( us03_n742 ) , .A1( us03_n784 ) );
  NOR2_X1 us03_U249 (.ZN( us03_n552 ) , .A1( us03_n784 ) , .A2( us03_n811 ) );
  NOR4_X1 us03_U25 (.A3( us03_n519 ) , .A1( us03_n520 ) , .ZN( us03_n521 ) , .A2( us03_n671 ) , .A4( us03_n767 ) );
  NOR2_X1 us03_U250 (.ZN( us03_n515 ) , .A1( us03_n706 ) , .A2( us03_n801 ) );
  NOR2_X1 us03_U251 (.ZN( us03_n556 ) , .A1( us03_n706 ) , .A2( us03_n814 ) );
  NOR2_X1 us03_U252 (.ZN( us03_n519 ) , .A1( us03_n788 ) , .A2( us03_n810 ) );
  INV_X1 us03_U253 (.A( us03_n803 ) , .ZN( us03_n858 ) );
  NOR2_X1 us03_U254 (.ZN( us03_n628 ) , .A1( us03_n745 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U255 (.ZN( us03_n713 ) , .A1( us03_n803 ) , .A2( us03_n815 ) );
  AOI21_X1 us03_U256 (.ZN( us03_n569 ) , .B2( us03_n695 ) , .B1( us03_n804 ) , .A( us03_n810 ) );
  NOR2_X1 us03_U257 (.ZN( us03_n653 ) , .A1( us03_n788 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U258 (.ZN( us03_n666 ) , .A2( us03_n706 ) , .A1( us03_n788 ) );
  NOR2_X1 us03_U259 (.ZN( us03_n654 ) , .A1( us03_n745 ) , .A2( us03_n778 ) );
  AOI222_X1 us03_U26 (.B2( us03_n636 ) , .ZN( us03_n642 ) , .B1( us03_n839 ) , .A1( us03_n840 ) , .C2( us03_n844 ) , .C1( us03_n861 ) , .A2( us03_n863 ) );
  NOR2_X1 us03_U260 (.ZN( us03_n554 ) , .A1( us03_n760 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U261 (.ZN( us03_n540 ) , .A1( us03_n760 ) , .A2( us03_n789 ) );
  NOR2_X1 us03_U262 (.ZN( us03_n699 ) , .A2( us03_n784 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U263 (.ZN( us03_n607 ) , .A2( us03_n722 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U264 (.A1( us03_n728 ) , .ZN( us03_n763 ) , .A2( us03_n784 ) );
  AOI21_X1 us03_U265 (.A( us03_n813 ) , .B2( us03_n814 ) , .B1( us03_n815 ) , .ZN( us03_n816 ) );
  NOR2_X1 us03_U266 (.ZN( us03_n577 ) , .A2( us03_n706 ) , .A1( us03_n728 ) );
  NOR2_X1 us03_U267 (.ZN( us03_n531 ) , .A2( us03_n722 ) , .A1( us03_n728 ) );
  AOI21_X1 us03_U268 (.B1( us03_n623 ) , .ZN( us03_n625 ) , .A( us03_n761 ) , .B2( us03_n812 ) );
  AOI21_X1 us03_U269 (.A( us03_n810 ) , .B2( us03_n811 ) , .B1( us03_n812 ) , .ZN( us03_n817 ) );
  NOR4_X1 us03_U27 (.A4( us03_n637 ) , .A3( us03_n638 ) , .A2( us03_n639 ) , .A1( us03_n640 ) , .ZN( us03_n641 ) );
  AOI21_X1 us03_U270 (.ZN( us03_n513 ) , .A( us03_n727 ) , .B1( us03_n748 ) , .B2( us03_n801 ) );
  AOI21_X1 us03_U271 (.ZN( us03_n497 ) , .B1( us03_n678 ) , .A( us03_n810 ) , .B2( us03_n814 ) );
  AOI21_X1 us03_U272 (.ZN( us03_n476 ) , .B2( us03_n695 ) , .A( us03_n747 ) , .B1( us03_n777 ) );
  NOR2_X1 us03_U273 (.ZN( us03_n580 ) , .A1( us03_n742 ) , .A2( us03_n813 ) );
  NOR2_X1 us03_U274 (.ZN( us03_n640 ) , .A2( us03_n786 ) , .A1( us03_n789 ) );
  AOI21_X1 us03_U275 (.ZN( us03_n591 ) , .B1( us03_n748 ) , .A( us03_n790 ) , .B2( us03_n811 ) );
  NOR2_X1 us03_U276 (.A2( us03_n706 ) , .A1( us03_n760 ) , .ZN( us03_n792 ) );
  AOI21_X1 us03_U277 (.ZN( us03_n624 ) , .B2( us03_n667 ) , .A( us03_n788 ) , .B1( us03_n789 ) );
  NOR2_X1 us03_U278 (.ZN( us03_n668 ) , .A1( us03_n788 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U279 (.ZN( us03_n518 ) , .A2( us03_n706 ) , .A1( us03_n812 ) );
  NOR3_X1 us03_U28 (.A2( us03_n605 ) , .A1( us03_n606 ) , .ZN( us03_n644 ) , .A3( us03_n720 ) );
  AOI21_X1 us03_U280 (.ZN( us03_n475 ) , .A( us03_n667 ) , .B1( us03_n748 ) , .B2( us03_n804 ) );
  NOR2_X1 us03_U281 (.ZN( us03_n557 ) , .A2( us03_n789 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U282 (.ZN( us03_n517 ) , .A2( us03_n697 ) , .A1( us03_n814 ) );
  NOR2_X1 us03_U283 (.ZN( us03_n681 ) , .A2( us03_n697 ) , .A1( us03_n801 ) );
  NOR2_X1 us03_U284 (.ZN( us03_n651 ) , .A1( us03_n760 ) , .A2( us03_n784 ) );
  INV_X1 us03_U285 (.A( us03_n811 ) , .ZN( us03_n834 ) );
  AOI21_X1 us03_U286 (.ZN( us03_n508 ) , .B2( us03_n667 ) , .A( us03_n728 ) , .B1( us03_n813 ) );
  AOI21_X1 us03_U287 (.ZN( us03_n537 ) , .B2( us03_n810 ) , .A( us03_n812 ) , .B1( us03_n813 ) );
  INV_X1 us03_U288 (.A( us03_n761 ) , .ZN( us03_n864 ) );
  AOI21_X1 us03_U289 (.ZN( us03_n538 ) , .A( us03_n761 ) , .B2( us03_n777 ) , .B1( us03_n815 ) );
  AOI221_X1 us03_U29 (.A( us03_n779 ) , .ZN( us03_n796 ) , .C2( us03_n835 ) , .B2( us03_n836 ) , .B1( us03_n863 ) , .C1( us03_n864 ) );
  NOR2_X1 us03_U290 (.ZN( us03_n579 ) , .A1( us03_n667 ) , .A2( us03_n786 ) );
  AOI21_X1 us03_U291 (.ZN( us03_n587 ) , .B2( us03_n697 ) , .B1( us03_n813 ) , .A( us03_n815 ) );
  AOI21_X1 us03_U292 (.B1( us03_n697 ) , .ZN( us03_n698 ) , .A( us03_n730 ) , .B2( us03_n761 ) );
  AOI21_X1 us03_U293 (.ZN( us03_n589 ) , .B2( us03_n761 ) , .A( us03_n783 ) , .B1( us03_n810 ) );
  AOI21_X1 us03_U294 (.ZN( us03_n496 ) , .A( us03_n722 ) , .B2( us03_n760 ) , .B1( us03_n812 ) );
  AOI21_X1 us03_U295 (.ZN( us03_n550 ) , .B1( us03_n667 ) , .A( us03_n695 ) , .B2( us03_n803 ) );
  NOR2_X1 us03_U296 (.ZN( us03_n545 ) , .A1( us03_n697 ) , .A2( us03_n742 ) );
  INV_X1 us03_U297 (.A( us03_n727 ) , .ZN( us03_n866 ) );
  INV_X1 us03_U298 (.A( us03_n789 ) , .ZN( us03_n871 ) );
  INV_X1 us03_U299 (.A( us03_n810 ) , .ZN( us03_n852 ) );
  NOR3_X1 us03_U3 (.ZN( us03_n596 ) , .A1( us03_n606 ) , .A3( us03_n721 ) , .A2( us03_n740 ) );
  NOR4_X1 us03_U30 (.A4( us03_n791 ) , .A3( us03_n792 ) , .A2( us03_n793 ) , .A1( us03_n794 ) , .ZN( us03_n795 ) );
  AOI21_X1 us03_U300 (.ZN( us03_n638 ) , .B2( us03_n745 ) , .A( us03_n790 ) , .B1( us03_n801 ) );
  AOI21_X1 us03_U301 (.ZN( us03_n647 ) , .B1( us03_n727 ) , .B2( us03_n761 ) , .A( us03_n811 ) );
  INV_X1 us03_U302 (.A( us03_n784 ) , .ZN( us03_n860 ) );
  NOR2_X1 us03_U303 (.ZN( us03_n683 ) , .A1( us03_n727 ) , .A2( us03_n814 ) );
  AOI21_X1 us03_U304 (.B1( us03_n684 ) , .ZN( us03_n685 ) , .A( us03_n726 ) , .B2( us03_n759 ) );
  AOI21_X1 us03_U305 (.ZN( us03_n567 ) , .B1( us03_n748 ) , .B2( us03_n760 ) , .A( us03_n778 ) );
  AOI21_X1 us03_U306 (.ZN( us03_n498 ) , .A( us03_n695 ) , .B1( us03_n706 ) , .B2( us03_n784 ) );
  NOR2_X1 us03_U307 (.ZN( us03_n566 ) , .A1( us03_n727 ) , .A2( us03_n760 ) );
  AOI21_X1 us03_U308 (.ZN( us03_n637 ) , .B2( us03_n747 ) , .A( us03_n786 ) , .B1( us03_n810 ) );
  NOR2_X1 us03_U309 (.ZN( us03_n564 ) , .A2( us03_n695 ) , .A1( us03_n761 ) );
  NOR4_X1 us03_U31 (.A4( us03_n774 ) , .A3( us03_n775 ) , .A1( us03_n776 ) , .ZN( us03_n797 ) , .A2( us03_n799 ) );
  NOR2_X1 us03_U310 (.ZN( us03_n578 ) , .A2( us03_n695 ) , .A1( us03_n789 ) );
  AOI21_X1 us03_U311 (.ZN( us03_n512 ) , .A( us03_n777 ) , .B2( us03_n790 ) , .B1( us03_n810 ) );
  INV_X1 us03_U312 (.A( us03_n697 ) , .ZN( us03_n851 ) );
  NOR2_X1 us03_U313 (.ZN( us03_n663 ) , .A1( us03_n778 ) , .A2( us03_n811 ) );
  AOI21_X1 us03_U314 (.ZN( us03_n448 ) , .B2( us03_n790 ) , .A( us03_n801 ) , .B1( us03_n813 ) );
  NOR2_X1 us03_U315 (.ZN( us03_n630 ) , .A2( us03_n695 ) , .A1( us03_n722 ) );
  AOI21_X1 us03_U316 (.ZN( us03_n562 ) , .B1( us03_n722 ) , .A( us03_n777 ) , .B2( us03_n789 ) );
  AOI21_X1 us03_U317 (.ZN( us03_n687 ) , .B2( us03_n747 ) , .B1( us03_n761 ) , .A( us03_n804 ) );
  NOR2_X1 us03_U318 (.ZN( us03_n527 ) , .A1( us03_n706 ) , .A2( us03_n777 ) );
  NOR2_X1 us03_U319 (.ZN( us03_n576 ) , .A1( us03_n706 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U32 (.ZN( us03_n802 ) , .A1( us03_n852 ) , .A2( us03_n859 ) );
  AOI21_X1 us03_U320 (.ZN( us03_n648 ) , .A( us03_n777 ) , .B1( us03_n790 ) , .B2( us03_n803 ) );
  NOR2_X1 us03_U321 (.ZN( us03_n682 ) , .A1( us03_n789 ) , .A2( us03_n811 ) );
  NOR2_X1 us03_U322 (.A2( us03_n811 ) , .A1( us03_n813 ) , .ZN( us03_n819 ) );
  AOI21_X1 us03_U323 (.A( us03_n788 ) , .B2( us03_n789 ) , .B1( us03_n790 ) , .ZN( us03_n791 ) );
  AOI21_X1 us03_U324 (.A( us03_n731 ) , .ZN( us03_n732 ) , .B2( us03_n778 ) , .B1( us03_n790 ) );
  NOR2_X1 us03_U325 (.ZN( us03_n565 ) , .A1( us03_n745 ) , .A2( us03_n803 ) );
  NOR2_X1 us03_U326 (.ZN( us03_n581 ) , .A1( us03_n790 ) , .A2( us03_n815 ) );
  NOR2_X1 us03_U327 (.ZN( us03_n532 ) , .A1( us03_n722 ) , .A2( us03_n786 ) );
  AOI21_X1 us03_U328 (.ZN( us03_n639 ) , .B1( us03_n678 ) , .A( us03_n789 ) , .B2( us03_n815 ) );
  NOR2_X1 us03_U329 (.ZN( us03_n709 ) , .A1( us03_n760 ) , .A2( us03_n761 ) );
  NAND4_X1 us03_U33 (.ZN( sa03_sr_7 ) , .A4( us03_n820 ) , .A3( us03_n821 ) , .A2( us03_n822 ) , .A1( us03_n823 ) );
  NOR2_X1 us03_U330 (.ZN( us03_n680 ) , .A2( us03_n706 ) , .A1( us03_n815 ) );
  INV_X1 us03_U331 (.A( us03_n695 ) , .ZN( us03_n836 ) );
  INV_X1 us03_U332 (.A( us03_n813 ) , .ZN( us03_n853 ) );
  AOI21_X1 us03_U333 (.ZN( us03_n440 ) , .A( us03_n697 ) , .B1( us03_n731 ) , .B2( us03_n748 ) );
  OAI21_X1 us03_U334 (.A( us03_n696 ) , .ZN( us03_n700 ) , .B2( us03_n748 ) , .B1( us03_n802 ) );
  OAI21_X1 us03_U335 (.ZN( us03_n696 ) , .B2( us03_n831 ) , .B1( us03_n836 ) , .A( us03_n858 ) );
  INV_X1 us03_U336 (.A( us03_n778 ) , .ZN( us03_n848 ) );
  AOI22_X1 us03_U337 (.A2( us03_n780 ) , .ZN( us03_n781 ) , .B2( us03_n829 ) , .A1( us03_n832 ) , .B1( us03_n861 ) );
  NAND2_X1 us03_U338 (.ZN( us03_n712 ) , .A1( us03_n726 ) , .A2( us03_n778 ) );
  NAND2_X1 us03_U339 (.ZN( us03_n751 ) , .A1( us03_n761 ) , .A2( us03_n803 ) );
  NOR4_X1 us03_U34 (.A4( us03_n816 ) , .A3( us03_n817 ) , .A2( us03_n818 ) , .A1( us03_n819 ) , .ZN( us03_n820 ) );
  NAND2_X1 us03_U340 (.A2( us03_n760 ) , .A1( us03_n804 ) , .ZN( us03_n808 ) );
  AOI21_X1 us03_U341 (.ZN( us03_n441 ) , .B1( us03_n787 ) , .B2( us03_n789 ) , .A( us03_n812 ) );
  OAI21_X1 us03_U343 (.A( us03_n785 ) , .B2( us03_n786 ) , .B1( us03_n787 ) , .ZN( us03_n793 ) );
  OAI21_X1 us03_U344 (.ZN( us03_n785 ) , .A( us03_n837 ) , .B1( us03_n861 ) , .B2( us03_n871 ) );
  AOI21_X1 us03_U345 (.ZN( us03_n495 ) , .A( us03_n777 ) , .B2( us03_n789 ) , .B1( us03_n802 ) );
  NAND2_X2 us03_U346 (.A2( us03_n439 ) , .A1( us03_n445 ) , .ZN( us03_n782 ) );
  INV_X1 us03_U347 (.A( us03_n783 ) , .ZN( us03_n844 ) );
  NOR2_X1 us03_U348 (.ZN( us03_n468 ) , .A2( us03_n777 ) , .A1( us03_n813 ) );
  OAI21_X1 us03_U349 (.A( us03_n729 ) , .B1( us03_n730 ) , .ZN( us03_n734 ) , .B2( us03_n803 ) );
  AOI222_X1 us03_U35 (.C2( us03_n807 ) , .B2( us03_n808 ) , .A2( us03_n809 ) , .ZN( us03_n821 ) , .C1( us03_n830 ) , .A1( us03_n837 ) , .B1( us03_n851 ) );
  OAI21_X1 us03_U350 (.ZN( us03_n729 ) , .A( us03_n831 ) , .B2( us03_n850 ) , .B1( us03_n871 ) );
  NOR2_X1 us03_U351 (.ZN( us03_n524 ) , .A1( us03_n722 ) , .A2( us03_n748 ) );
  NOR2_X1 us03_U352 (.ZN( us03_n710 ) , .A2( us03_n722 ) , .A1( us03_n788 ) );
  NOR2_X1 us03_U353 (.ZN( us03_n482 ) , .A1( us03_n786 ) , .A2( us03_n803 ) );
  NAND2_X1 us03_U354 (.A1( us03_n697 ) , .A2( us03_n727 ) , .ZN( us03_n780 ) );
  NOR2_X1 us03_U355 (.ZN( us03_n516 ) , .A1( us03_n706 ) , .A2( us03_n786 ) );
  NAND2_X1 us03_U356 (.ZN( us03_n669 ) , .A1( us03_n804 ) , .A2( us03_n814 ) );
  NAND2_X1 us03_U357 (.A2( us03_n747 ) , .A1( us03_n784 ) , .ZN( us03_n807 ) );
  INV_X1 us03_U358 (.A( us03_n722 ) , .ZN( us03_n854 ) );
  INV_X1 us03_U359 (.A( us03_n815 ) , .ZN( us03_n842 ) );
  AOI211_X1 us03_U36 (.B( us03_n805 ) , .A( us03_n806 ) , .ZN( us03_n822 ) , .C1( us03_n840 ) , .C2( us03_n848 ) );
  AND2_X1 us03_U360 (.ZN( us03_n730 ) , .A1( us03_n777 ) , .A2( us03_n783 ) );
  NAND2_X1 us03_U366 (.A1( us03_n450 ) , .A2( us03_n463 ) , .ZN( us03_n667 ) );
  NOR2_X1 us03_U37 (.ZN( us03_n746 ) , .A1( us03_n859 ) , .A2( us03_n860 ) );
  NAND2_X1 us03_U372 (.A2( us03_n462 ) , .A1( us03_n463 ) , .ZN( us03_n810 ) );
  NAND2_X1 us03_U373 (.A1( us03_n439 ) , .A2( us03_n458 ) , .ZN( us03_n697 ) );
  NOR2_X1 us03_U38 (.ZN( us03_n623 ) , .A2( us03_n834 ) , .A1( us03_n837 ) );
  NAND2_X2 us03_U385 (.A2( us03_n439 ) , .A1( us03_n450 ) , .ZN( us03_n789 ) );
  NAND2_X2 us03_U388 (.A1( us03_n439 ) , .A2( us03_n462 ) , .ZN( us03_n706 ) );
  NAND4_X1 us03_U39 (.A4( us03_n601 ) , .A3( us03_n602 ) , .A2( us03_n603 ) , .A1( us03_n604 ) , .ZN( us03_n720 ) );
  NAND2_X2 us03_U390 (.A2( us03_n458 ) , .A1( us03_n463 ) , .ZN( us03_n778 ) );
  NOR2_X1 us03_U397 (.A2( sa03_4 ) , .A1( sa03_5 ) , .ZN( us03_n439 ) );
  NOR3_X1 us03_U4 (.A3( us03_n798 ) , .A2( us03_n799 ) , .A1( us03_n800 ) , .ZN( us03_n823 ) );
  NOR3_X1 us03_U40 (.A1( us03_n597 ) , .ZN( us03_n602 ) , .A3( us03_n661 ) , .A2( us03_n768 ) );
  NOR4_X1 us03_U41 (.A3( us03_n598 ) , .A2( us03_n599 ) , .A1( us03_n600 ) , .ZN( us03_n601 ) , .A4( us03_n653 ) );
  AOI222_X1 us03_U412 (.ZN( us03_n603 ) , .B2( us03_n669 ) , .B1( us03_n751 ) , .C2( us03_n829 ) , .A1( us03_n831 ) , .A2( us03_n860 ) , .C1( us03_n861 ) );
  AOI222_X1 us03_U413 (.ZN( us03_n511 ) , .C1( us03_n830 ) , .B2( us03_n835 ) , .A2( us03_n841 ) , .C2( us03_n860 ) , .B1( us03_n861 ) , .A1( us03_n864 ) );
  AOI221_X1 us03_U414 (.A( us03_n481 ) , .ZN( us03_n486 ) , .B1( us03_n829 ) , .C2( us03_n842 ) , .C1( us03_n850 ) , .B2( us03_n860 ) );
  NOR2_X1 us03_U415 (.ZN( us03_n787 ) , .A2( us03_n860 ) , .A1( us03_n866 ) );
  NAND4_X1 us03_U416 (.ZN( sa03_sr_2 ) , .A4( us03_n641 ) , .A3( us03_n642 ) , .A2( us03_n643 ) , .A1( us03_n644 ) );
  OAI221_X1 us03_U417 (.A( us03_n781 ) , .C2( us03_n782 ) , .B2( us03_n783 ) , .B1( us03_n784 ) , .ZN( us03_n794 ) , .C1( us03_n811 ) );
  NAND2_X1 us03_U418 (.A1( us03_n727 ) , .A2( us03_n782 ) , .ZN( us03_n809 ) );
  OAI22_X1 us03_U419 (.ZN( us03_n586 ) , .A2( us03_n745 ) , .B2( us03_n760 ) , .A1( us03_n761 ) , .B1( us03_n782 ) );
  AOI222_X1 us03_U42 (.ZN( us03_n604 ) , .A1( us03_n828 ) , .C2( us03_n835 ) , .B1( us03_n840 ) , .A2( us03_n854 ) , .B2( us03_n859 ) , .C1( us03_n866 ) );
  OAI221_X1 us03_U420 (.A( us03_n694 ) , .ZN( us03_n701 ) , .C2( us03_n782 ) , .C1( us03_n783 ) , .B1( us03_n784 ) , .B2( us03_n804 ) );
  AOI21_X1 us03_U421 (.ZN( us03_n590 ) , .B1( us03_n726 ) , .B2( us03_n782 ) , .A( us03_n788 ) );
  AOI21_X1 us03_U422 (.ZN( us03_n621 ) , .B1( us03_n697 ) , .A( us03_n777 ) , .B2( us03_n782 ) );
  AOI21_X1 us03_U423 (.ZN( us03_n646 ) , .A( us03_n760 ) , .B2( us03_n782 ) , .B1( us03_n790 ) );
  OAI22_X1 us03_U424 (.ZN( us03_n679 ) , .A1( us03_n697 ) , .A2( us03_n728 ) , .B2( us03_n782 ) , .B1( us03_n815 ) );
  OAI21_X1 us03_U425 (.A( us03_n611 ) , .ZN( us03_n614 ) , .B1( us03_n623 ) , .B2( us03_n782 ) );
  NOR2_X1 us03_U426 (.ZN( us03_n608 ) , .A1( us03_n782 ) , .A2( us03_n814 ) );
  OAI222_X1 us03_U427 (.A2( us03_n667 ) , .ZN( us03_n672 ) , .B1( us03_n745 ) , .B2( us03_n782 ) , .C2( us03_n786 ) , .C1( us03_n813 ) , .A1( us03_n815 ) );
  NOR2_X1 us03_U428 (.ZN( us03_n649 ) , .A1( us03_n782 ) , .A2( us03_n786 ) );
  NOR2_X1 us03_U429 (.ZN( us03_n598 ) , .A2( us03_n695 ) , .A1( us03_n782 ) );
  NAND4_X1 us03_U43 (.ZN( sa03_sr_3 ) , .A4( us03_n702 ) , .A3( us03_n703 ) , .A2( us03_n704 ) , .A1( us03_n705 ) );
  NOR2_X1 us03_U430 (.ZN( us03_n551 ) , .A2( us03_n742 ) , .A1( us03_n782 ) );
  INV_X1 us03_U431 (.A( us03_n782 ) , .ZN( us03_n859 ) );
  AOI221_X1 us03_U432 (.A( us03_n574 ) , .ZN( us03_n585 ) , .B2( us03_n829 ) , .C2( us03_n841 ) , .B1( us03_n852 ) , .C1( us03_n859 ) );
  AOI21_X1 us03_U433 (.ZN( us03_n574 ) , .B2( us03_n722 ) , .B1( us03_n746 ) , .A( us03_n783 ) );
  AOI211_X1 us03_U434 (.A( us03_n635 ) , .ZN( us03_n643 ) , .B( us03_n741 ) , .C2( us03_n837 ) , .C1( us03_n852 ) );
  NAND4_X1 us03_U435 (.A4( us03_n631 ) , .A3( us03_n632 ) , .A2( us03_n633 ) , .A1( us03_n634 ) , .ZN( us03_n741 ) );
  NAND3_X1 us03_U437 (.ZN( sa03_sr_6 ) , .A3( us03_n795 ) , .A2( us03_n796 ) , .A1( us03_n797 ) );
  NAND3_X1 us03_U438 (.ZN( sa03_sr_5 ) , .A3( us03_n756 ) , .A2( us03_n757 ) , .A1( us03_n758 ) );
  NAND3_X1 us03_U439 (.ZN( sa03_sr_4 ) , .A3( us03_n736 ) , .A2( us03_n737 ) , .A1( us03_n738 ) );
  NOR4_X1 us03_U44 (.A4( us03_n698 ) , .A3( us03_n699 ) , .A2( us03_n700 ) , .A1( us03_n701 ) , .ZN( us03_n702 ) );
  NAND3_X1 us03_U440 (.A3( us03_n673 ) , .A2( us03_n674 ) , .A1( us03_n675 ) , .ZN( us03_n805 ) );
  NAND3_X1 us03_U441 (.ZN( us03_n636 ) , .A3( us03_n706 ) , .A2( us03_n722 ) , .A1( us03_n790 ) );
  NAND3_X1 us03_U442 (.A3( us03_n616 ) , .A2( us03_n617 ) , .A1( us03_n618 ) , .ZN( us03_n723 ) );
  NAND3_X1 us03_U443 (.A3( us03_n583 ) , .A2( us03_n584 ) , .A1( us03_n585 ) , .ZN( us03_n619 ) );
  NAND3_X1 us03_U444 (.ZN( us03_n563 ) , .A3( us03_n678 ) , .A2( us03_n748 ) , .A1( us03_n783 ) );
  NAND3_X1 us03_U445 (.A3( us03_n521 ) , .A2( us03_n522 ) , .A1( us03_n523 ) , .ZN( us03_n740 ) );
  NAND3_X1 us03_U446 (.A3( us03_n510 ) , .A1( us03_n511 ) , .ZN( us03_n606 ) , .A2( us03_n869 ) );
  NAND3_X1 us03_U447 (.A3( us03_n465 ) , .A2( us03_n466 ) , .A1( us03_n467 ) , .ZN( us03_n775 ) );
  AOI211_X1 us03_U45 (.B( us03_n692 ) , .A( us03_n693 ) , .ZN( us03_n703 ) , .C2( us03_n829 ) , .C1( us03_n849 ) );
  NOR2_X1 us03_U46 (.ZN( us03_n705 ) , .A2( us03_n774 ) , .A1( us03_n798 ) );
  AOI222_X1 us03_U47 (.ZN( us03_n467 ) , .B1( us03_n830 ) , .A1( us03_n837 ) , .C1( us03_n840 ) , .C2( us03_n849 ) , .A2( us03_n853 ) , .B2( us03_n863 ) );
  NOR4_X1 us03_U48 (.A1( us03_n464 ) , .ZN( us03_n465 ) , .A4( us03_n540 ) , .A2( us03_n552 ) , .A3( us03_n612 ) );
  AOI221_X1 us03_U49 (.ZN( us03_n466 ) , .C2( us03_n712 ) , .B2( us03_n829 ) , .C1( us03_n843 ) , .B1( us03_n858 ) , .A( us03_n862 ) );
  NOR3_X1 us03_U5 (.ZN( us03_n502 ) , .A2( us03_n677 ) , .A3( us03_n775 ) , .A1( us03_n874 ) );
  NOR4_X1 us03_U50 (.A4( us03_n575 ) , .A3( us03_n576 ) , .A2( us03_n577 ) , .ZN( us03_n584 ) , .A1( us03_n681 ) );
  NOR4_X1 us03_U51 (.A1( us03_n582 ) , .ZN( us03_n583 ) , .A3( us03_n650 ) , .A2( us03_n660 ) , .A4( us03_n765 ) );
  NAND4_X1 us03_U52 (.A4( us03_n483 ) , .A3( us03_n484 ) , .A2( us03_n485 ) , .A1( us03_n486 ) , .ZN( us03_n776 ) );
  NOR4_X1 us03_U53 (.A4( us03_n482 ) , .ZN( us03_n485 ) , .A1( us03_n564 ) , .A2( us03_n579 ) , .A3( us03_n600 ) );
  NOR4_X1 us03_U54 (.ZN( us03_n484 ) , .A1( us03_n505 ) , .A2( us03_n517 ) , .A4( us03_n544 ) , .A3( us03_n609 ) );
  NOR4_X1 us03_U55 (.ZN( us03_n483 ) , .A2( us03_n531 ) , .A1( us03_n556 ) , .A3( us03_n629 ) , .A4( us03_n716 ) );
  AOI211_X1 us03_U56 (.B( us03_n621 ) , .A( us03_n622 ) , .ZN( us03_n633 ) , .C2( us03_n834 ) , .C1( us03_n861 ) );
  NOR4_X1 us03_U57 (.A4( us03_n627 ) , .A3( us03_n628 ) , .A2( us03_n629 ) , .A1( us03_n630 ) , .ZN( us03_n631 ) );
  NOR4_X1 us03_U58 (.A4( us03_n624 ) , .A3( us03_n625 ) , .A2( us03_n626 ) , .ZN( us03_n632 ) , .A1( us03_n662 ) );
  NAND4_X1 us03_U59 (.A4( us03_n655 ) , .A3( us03_n656 ) , .A2( us03_n657 ) , .A1( us03_n658 ) , .ZN( us03_n798 ) );
  INV_X1 us03_U6 (.A( us03_n704 ) , .ZN( us03_n874 ) );
  NOR3_X1 us03_U60 (.A3( us03_n646 ) , .A2( us03_n647 ) , .A1( us03_n648 ) , .ZN( us03_n657 ) );
  NOR3_X1 us03_U61 (.A3( us03_n649 ) , .A2( us03_n650 ) , .A1( us03_n651 ) , .ZN( us03_n656 ) );
  NOR3_X1 us03_U62 (.A3( us03_n652 ) , .A2( us03_n653 ) , .A1( us03_n654 ) , .ZN( us03_n655 ) );
  NAND4_X1 us03_U63 (.A4( us03_n558 ) , .A3( us03_n559 ) , .A2( us03_n560 ) , .A1( us03_n561 ) , .ZN( us03_n605 ) );
  NOR4_X1 us03_U64 (.A4( us03_n554 ) , .A3( us03_n555 ) , .A2( us03_n556 ) , .A1( us03_n557 ) , .ZN( us03_n558 ) );
  NOR4_X1 us03_U65 (.ZN( us03_n559 ) , .A1( us03_n651 ) , .A3( us03_n659 ) , .A4( us03_n683 ) , .A2( us03_n766 ) );
  NOR4_X1 us03_U66 (.A4( us03_n550 ) , .A3( us03_n551 ) , .A2( us03_n552 ) , .A1( us03_n553 ) , .ZN( us03_n560 ) );
  NAND4_X1 us03_U67 (.A4( us03_n770 ) , .A3( us03_n771 ) , .A2( us03_n772 ) , .A1( us03_n773 ) , .ZN( us03_n799 ) );
  NOR3_X1 us03_U68 (.A3( us03_n763 ) , .A2( us03_n764 ) , .A1( us03_n765 ) , .ZN( us03_n771 ) );
  NOR4_X1 us03_U69 (.A4( us03_n766 ) , .A3( us03_n767 ) , .A2( us03_n768 ) , .A1( us03_n769 ) , .ZN( us03_n770 ) );
  NOR3_X1 us03_U7 (.A3( us03_n619 ) , .A2( us03_n620 ) , .ZN( us03_n634 ) , .A1( us03_n723 ) );
  AOI222_X1 us03_U70 (.ZN( us03_n773 ) , .A1( us03_n828 ) , .C1( us03_n832 ) , .B2( us03_n839 ) , .A2( us03_n848 ) , .B1( us03_n859 ) , .C2( us03_n871 ) );
  NOR4_X1 us03_U71 (.A4( us03_n507 ) , .A2( us03_n508 ) , .A1( us03_n509 ) , .ZN( us03_n510 ) , .A3( us03_n668 ) );
  INV_X1 us03_U72 (.A( us03_n503 ) , .ZN( us03_n869 ) );
  NOR4_X1 us03_U73 (.A4( us03_n663 ) , .A3( us03_n664 ) , .A2( us03_n665 ) , .A1( us03_n666 ) , .ZN( us03_n674 ) );
  NOR4_X1 us03_U74 (.A4( us03_n659 ) , .A3( us03_n660 ) , .A2( us03_n661 ) , .A1( us03_n662 ) , .ZN( us03_n675 ) );
  NOR4_X1 us03_U75 (.A3( us03_n671 ) , .A1( us03_n672 ) , .ZN( us03_n673 ) , .A4( us03_n713 ) , .A2( us03_n857 ) );
  NOR2_X1 us03_U76 (.ZN( us03_n759 ) , .A1( us03_n831 ) , .A2( us03_n832 ) );
  NOR4_X1 us03_U77 (.A4( us03_n732 ) , .A3( us03_n733 ) , .A2( us03_n734 ) , .A1( us03_n735 ) , .ZN( us03_n736 ) );
  AOI211_X1 us03_U78 (.B( us03_n723 ) , .A( us03_n724 ) , .ZN( us03_n737 ) , .C1( us03_n841 ) , .C2( us03_n853 ) );
  NOR3_X1 us03_U79 (.A3( us03_n720 ) , .A1( us03_n721 ) , .ZN( us03_n738 ) , .A2( us03_n739 ) );
  NOR2_X1 us03_U8 (.ZN( us03_n573 ) , .A1( us03_n620 ) , .A2( us03_n743 ) );
  NOR4_X1 us03_U80 (.A3( us03_n753 ) , .A2( us03_n754 ) , .A1( us03_n755 ) , .ZN( us03_n756 ) , .A4( us03_n867 ) );
  AOI211_X1 us03_U81 (.B( us03_n743 ) , .A( us03_n744 ) , .ZN( us03_n757 ) , .C1( us03_n830 ) , .C2( us03_n851 ) );
  NOR3_X1 us03_U82 (.A3( us03_n739 ) , .A2( us03_n740 ) , .A1( us03_n741 ) , .ZN( us03_n758 ) );
  NAND4_X1 us03_U83 (.A4( us03_n454 ) , .A3( us03_n455 ) , .A2( us03_n456 ) , .A1( us03_n457 ) , .ZN( us03_n677 ) );
  NOR3_X1 us03_U84 (.ZN( us03_n455 ) , .A3( us03_n528 ) , .A1( us03_n553 ) , .A2( us03_n568 ) );
  AOI221_X1 us03_U85 (.A( us03_n448 ) , .ZN( us03_n457 ) , .C2( us03_n751 ) , .B1( us03_n830 ) , .C1( us03_n840 ) , .B2( us03_n859 ) );
  NOR4_X1 us03_U86 (.ZN( us03_n456 ) , .A2( us03_n507 ) , .A1( us03_n597 ) , .A4( us03_n626 ) , .A3( us03_n709 ) );
  NAND4_X1 us03_U87 (.A4( us03_n533 ) , .A3( us03_n534 ) , .A2( us03_n535 ) , .A1( us03_n536 ) , .ZN( us03_n620 ) );
  NOR4_X1 us03_U88 (.A4( us03_n524 ) , .A2( us03_n525 ) , .A1( us03_n526 ) , .ZN( us03_n536 ) , .A3( us03_n699 ) );
  NOR4_X1 us03_U89 (.A1( us03_n529 ) , .ZN( us03_n534 ) , .A2( us03_n652 ) , .A4( us03_n666 ) , .A3( us03_n763 ) );
  NOR2_X1 us03_U9 (.A1( us03_n676 ) , .ZN( us03_n691 ) , .A2( us03_n805 ) );
  NOR4_X1 us03_U90 (.A4( us03_n527 ) , .A3( us03_n528 ) , .ZN( us03_n535 ) , .A2( us03_n682 ) , .A1( us03_n792 ) );
  NAND4_X1 us03_U91 (.A4( us03_n477 ) , .A3( us03_n478 ) , .A2( us03_n479 ) , .A1( us03_n480 ) , .ZN( us03_n692 ) );
  NOR3_X1 us03_U92 (.ZN( us03_n478 ) , .A2( us03_n506 ) , .A3( us03_n599 ) , .A1( us03_n608 ) );
  AOI211_X1 us03_U93 (.B( us03_n475 ) , .A( us03_n476 ) , .ZN( us03_n480 ) , .C2( us03_n831 ) , .C1( us03_n859 ) );
  NOR4_X1 us03_U94 (.ZN( us03_n479 ) , .A3( us03_n530 ) , .A4( us03_n543 ) , .A2( us03_n565 ) , .A1( us03_n715 ) );
  NAND4_X1 us03_U95 (.A4( us03_n546 ) , .A3( us03_n547 ) , .A2( us03_n548 ) , .A1( us03_n549 ) , .ZN( us03_n743 ) );
  NOR3_X1 us03_U96 (.ZN( us03_n547 ) , .A2( us03_n649 ) , .A1( us03_n665 ) , .A3( us03_n769 ) );
  AOI211_X1 us03_U97 (.B( us03_n537 ) , .A( us03_n538 ) , .ZN( us03_n549 ) , .C2( us03_n837 ) , .C1( us03_n849 ) );
  NOR4_X1 us03_U98 (.A4( us03_n542 ) , .A3( us03_n543 ) , .A2( us03_n544 ) , .A1( us03_n545 ) , .ZN( us03_n546 ) );
  NOR4_X1 us03_U99 (.ZN( us03_n618 ) , .A1( us03_n654 ) , .A3( us03_n664 ) , .A4( us03_n680 ) , .A2( us03_n764 ) );
endmodule

